// (C) 1992-2014 Altera Corporation. All rights reserved.                         
// Your use of Altera Corporation's design tools, logic functions and other       
// software and tools, and its AMPP partner logic functions, and any output       
// files any of the foregoing (including device programming or simulation         
// files), and any associated documentation or information are expressly subject  
// to the terms and conditions of the Altera Program License Subscription         
// Agreement, Altera MegaCore Function License Agreement, or other applicable     
// license agreement, including, without limitation, that your use is for the     
// sole purpose of programming logic devices manufactured by Altera and sold by   
// Altera or its authorized distributors.  Please refer to the applicable         
// agreement for further details.                                                 
    

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

module Matmul_basic_block_0
	(
		input 		clock,
		input 		resetn,
		input 		start,
		input [31:0] 		input_c1f2,
		input 		valid_in,
		output 		stall_out,
		input [31:0] 		input_global_id_0,
		input [31:0] 		input_global_id_1,
		output 		valid_out,
		input 		stall_in,
		output 		lvb_bb0_cmp3,
		output 		lvb_bb0_cmp3_NEG,
		output [31:0] 		lvb_input_global_id_0,
		output [31:0] 		lvb_input_global_id_1,
		input [31:0] 		workgroup_size
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_global_id_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_global_id_0_staging_reg_NO_SHIFT_REG <= input_global_id_0;
				input_global_id_1_staging_reg_NO_SHIFT_REG <= input_global_id_1;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp3_inputs_ready;
 reg local_bb0_cmp3_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp3_valid_out_0_NO_SHIFT_REG;
wire local_bb0_cmp3_stall_in_0;
 reg local_bb0_cmp3_valid_out_1_NO_SHIFT_REG;
wire local_bb0_cmp3_stall_in_1;
wire local_bb0_cmp3_output_regs_ready;
 reg local_bb0_cmp3_NO_SHIFT_REG;
wire local_bb0_cmp3_causedstall;

assign local_bb0_cmp3_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb0_cmp3_output_regs_ready = (~(local_bb0_cmp3_wii_reg_NO_SHIFT_REG) & ((~(local_bb0_cmp3_valid_out_0_NO_SHIFT_REG) | ~(local_bb0_cmp3_stall_in_0)) & (~(local_bb0_cmp3_valid_out_1_NO_SHIFT_REG) | ~(local_bb0_cmp3_stall_in_1))));
assign merge_node_stall_in_0 = (~(local_bb0_cmp3_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp3_output_regs_ready) | ~(local_bb0_cmp3_inputs_ready)));
assign local_bb0_cmp3_causedstall = (local_bb0_cmp3_inputs_ready && (~(local_bb0_cmp3_output_regs_ready) && !(~(local_bb0_cmp3_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp3_NO_SHIFT_REG <= 'x;
		local_bb0_cmp3_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb0_cmp3_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp3_NO_SHIFT_REG <= 'x;
			local_bb0_cmp3_valid_out_0_NO_SHIFT_REG <= 1'b0;
			local_bb0_cmp3_valid_out_1_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp3_output_regs_ready)
			begin
				local_bb0_cmp3_NO_SHIFT_REG <= ($signed(input_c1f2) > $signed(32'h0));
				local_bb0_cmp3_valid_out_0_NO_SHIFT_REG <= local_bb0_cmp3_inputs_ready;
				local_bb0_cmp3_valid_out_1_NO_SHIFT_REG <= local_bb0_cmp3_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp3_stall_in_0))
				begin
					local_bb0_cmp3_valid_out_0_NO_SHIFT_REG <= local_bb0_cmp3_wii_reg_NO_SHIFT_REG;
				end
				if (~(local_bb0_cmp3_stall_in_1))
				begin
					local_bb0_cmp3_valid_out_1_NO_SHIFT_REG <= local_bb0_cmp3_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp3_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp3_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp3_inputs_ready)
			begin
				local_bb0_cmp3_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb0_cmp3_NEG_inputs_ready;
 reg local_bb0_cmp3_NEG_wii_reg_NO_SHIFT_REG;
 reg local_bb0_cmp3_NEG_valid_out_NO_SHIFT_REG;
wire local_bb0_cmp3_NEG_stall_in;
wire local_bb0_cmp3_NEG_output_regs_ready;
 reg local_bb0_cmp3_NEG_NO_SHIFT_REG;
wire local_bb0_cmp3_NEG_causedstall;

assign local_bb0_cmp3_NEG_inputs_ready = local_bb0_cmp3_valid_out_0_NO_SHIFT_REG;
assign local_bb0_cmp3_NEG_output_regs_ready = (~(local_bb0_cmp3_NEG_wii_reg_NO_SHIFT_REG) & (&(~(local_bb0_cmp3_NEG_valid_out_NO_SHIFT_REG) | ~(local_bb0_cmp3_NEG_stall_in))));
assign local_bb0_cmp3_stall_in_0 = (~(local_bb0_cmp3_NEG_wii_reg_NO_SHIFT_REG) & (~(local_bb0_cmp3_NEG_output_regs_ready) | ~(local_bb0_cmp3_NEG_inputs_ready)));
assign local_bb0_cmp3_NEG_causedstall = (local_bb0_cmp3_NEG_inputs_ready && (~(local_bb0_cmp3_NEG_output_regs_ready) && !(~(local_bb0_cmp3_NEG_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp3_NEG_NO_SHIFT_REG <= 'x;
		local_bb0_cmp3_NEG_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp3_NEG_NO_SHIFT_REG <= 'x;
			local_bb0_cmp3_NEG_valid_out_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp3_NEG_output_regs_ready)
			begin
				local_bb0_cmp3_NEG_NO_SHIFT_REG <= (local_bb0_cmp3_NO_SHIFT_REG ^ 1'b1);
				local_bb0_cmp3_NEG_valid_out_NO_SHIFT_REG <= local_bb0_cmp3_NEG_inputs_ready;
			end
			else
			begin
				if (~(local_bb0_cmp3_NEG_stall_in))
				begin
					local_bb0_cmp3_NEG_valid_out_NO_SHIFT_REG <= local_bb0_cmp3_NEG_wii_reg_NO_SHIFT_REG;
				end
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb0_cmp3_NEG_wii_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (start)
		begin
			local_bb0_cmp3_NEG_wii_reg_NO_SHIFT_REG <= 1'b0;
		end
		else
		begin
			if (local_bb0_cmp3_NEG_inputs_ready)
			begin
				local_bb0_cmp3_NEG_wii_reg_NO_SHIFT_REG <= 1'b1;
			end
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg lvb_bb0_cmp3_reg_NO_SHIFT_REG;
 reg lvb_bb0_cmp3_NEG_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_1_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb0_cmp3_NEG_valid_out_NO_SHIFT_REG & merge_node_valid_out_1_NO_SHIFT_REG & local_bb0_cmp3_valid_out_1_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb0_cmp3_NEG_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign merge_node_stall_in_1 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb0_cmp3_stall_in_1 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb0_cmp3 = lvb_bb0_cmp3_reg_NO_SHIFT_REG;
assign lvb_bb0_cmp3_NEG = lvb_bb0_cmp3_NEG_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0 = lvb_input_global_id_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1 = lvb_input_global_id_1_reg_NO_SHIFT_REG;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb0_cmp3_reg_NO_SHIFT_REG <= 'x;
		lvb_bb0_cmp3_NEG_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_1_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb0_cmp3_reg_NO_SHIFT_REG <= local_bb0_cmp3_NO_SHIFT_REG;
			lvb_bb0_cmp3_NEG_reg_NO_SHIFT_REG <= local_bb0_cmp3_NEG_NO_SHIFT_REG;
			lvb_input_global_id_0_reg_NO_SHIFT_REG <= local_lvm_input_global_id_0_NO_SHIFT_REG;
			lvb_input_global_id_1_reg_NO_SHIFT_REG <= local_lvm_input_global_id_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

module Matmul_basic_block_1
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_c1f2,
		input 		input_wii_cmp3,
		input 		input_wii_cmp3_NEG,
		input 		valid_in,
		output 		stall_out,
		input [31:0] 		input_global_id_0,
		input [31:0] 		input_global_id_1,
		output 		valid_out,
		input 		stall_in,
		output [63:0] 		lvb_bb1_var_,
		output [31:0] 		lvb_input_global_id_0,
		output [31:0] 		lvb_input_global_id_1,
		input [31:0] 		workgroup_size,
		input 		start
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_global_id_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_global_id_0_staging_reg_NO_SHIFT_REG <= input_global_id_0;
				input_global_id_1_staging_reg_NO_SHIFT_REG <= input_global_id_1;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements a registered operation.
// 
wire local_bb1_mul_inputs_ready;
 reg local_bb1_mul_valid_out_NO_SHIFT_REG;
wire local_bb1_mul_stall_in;
wire local_bb1_mul_output_regs_ready;
wire [31:0] local_bb1_mul;
 reg local_bb1_mul_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb1_mul_valid_pipe_1_NO_SHIFT_REG;
wire local_bb1_mul_causedstall;

acl_int_mult32s_s5 int_module_local_bb1_mul (
	.clock(clock),
	.dataa(local_lvm_input_global_id_1_NO_SHIFT_REG),
	.datab(input_c1f2),
	.enable(local_bb1_mul_output_regs_ready),
	.result(local_bb1_mul)
);

defparam int_module_local_bb1_mul.INPUT1_WIDTH = 32;
defparam int_module_local_bb1_mul.INPUT2_WIDTH = 32;

assign local_bb1_mul_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb1_mul_output_regs_ready = (&(~(local_bb1_mul_valid_out_NO_SHIFT_REG) | ~(local_bb1_mul_stall_in)));
assign merge_node_stall_in_0 = (~(local_bb1_mul_output_regs_ready) | ~(local_bb1_mul_inputs_ready));
assign local_bb1_mul_causedstall = (local_bb1_mul_inputs_ready && (~(local_bb1_mul_output_regs_ready) && !(~(local_bb1_mul_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_mul_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb1_mul_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_mul_output_regs_ready)
		begin
			local_bb1_mul_valid_pipe_0_NO_SHIFT_REG <= local_bb1_mul_inputs_ready;
			local_bb1_mul_valid_pipe_1_NO_SHIFT_REG <= local_bb1_mul_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb1_mul_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb1_mul_output_regs_ready)
		begin
			local_bb1_mul_valid_out_NO_SHIFT_REG <= local_bb1_mul_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb1_mul_stall_in))
			begin
				local_bb1_mul_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_input_global_id_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_1to4_input_global_id_0_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_input_global_id_0_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_input_global_id_0_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_lvm_input_global_id_0_NO_SHIFT_REG),
	.data_out(rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_1_NO_SHIFT_REG;
assign merge_node_stall_in_1 = rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_stall_in_reg_4_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_stall_in_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_valid_out_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_valid_out_reg_4_NO_SHIFT_REG;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_input_global_id_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_1_0_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_1_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_1_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_1_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_1_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_1_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_1to4_input_global_id_1_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_input_global_id_1_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_input_global_id_1_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_input_global_id_1_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_input_global_id_1_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_lvm_input_global_id_1_NO_SHIFT_REG),
	.data_out(rnode_1to4_input_global_id_1_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_input_global_id_1_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_input_global_id_1_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_1to4_input_global_id_1_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_input_global_id_1_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_input_global_id_1_0_reg_4_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_2_NO_SHIFT_REG;
assign merge_node_stall_in_2 = rnode_1to4_input_global_id_1_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_1_0_NO_SHIFT_REG = rnode_1to4_input_global_id_1_0_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_1_0_stall_in_reg_4_NO_SHIFT_REG = rnode_1to4_input_global_id_1_0_stall_in_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_1_0_valid_out_NO_SHIFT_REG = rnode_1to4_input_global_id_1_0_valid_out_reg_4_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb1_var__valid_out;
wire local_bb1_var__stall_in;
wire local_bb1_var__inputs_ready;
wire local_bb1_var__stall_local;
wire [63:0] local_bb1_var_;

assign local_bb1_var__inputs_ready = local_bb1_mul_valid_out_NO_SHIFT_REG;
assign local_bb1_var_[32] = local_bb1_mul[31];
assign local_bb1_var_[33] = local_bb1_mul[31];
assign local_bb1_var_[34] = local_bb1_mul[31];
assign local_bb1_var_[35] = local_bb1_mul[31];
assign local_bb1_var_[36] = local_bb1_mul[31];
assign local_bb1_var_[37] = local_bb1_mul[31];
assign local_bb1_var_[38] = local_bb1_mul[31];
assign local_bb1_var_[39] = local_bb1_mul[31];
assign local_bb1_var_[40] = local_bb1_mul[31];
assign local_bb1_var_[41] = local_bb1_mul[31];
assign local_bb1_var_[42] = local_bb1_mul[31];
assign local_bb1_var_[43] = local_bb1_mul[31];
assign local_bb1_var_[44] = local_bb1_mul[31];
assign local_bb1_var_[45] = local_bb1_mul[31];
assign local_bb1_var_[46] = local_bb1_mul[31];
assign local_bb1_var_[47] = local_bb1_mul[31];
assign local_bb1_var_[48] = local_bb1_mul[31];
assign local_bb1_var_[49] = local_bb1_mul[31];
assign local_bb1_var_[50] = local_bb1_mul[31];
assign local_bb1_var_[51] = local_bb1_mul[31];
assign local_bb1_var_[52] = local_bb1_mul[31];
assign local_bb1_var_[53] = local_bb1_mul[31];
assign local_bb1_var_[54] = local_bb1_mul[31];
assign local_bb1_var_[55] = local_bb1_mul[31];
assign local_bb1_var_[56] = local_bb1_mul[31];
assign local_bb1_var_[57] = local_bb1_mul[31];
assign local_bb1_var_[58] = local_bb1_mul[31];
assign local_bb1_var_[59] = local_bb1_mul[31];
assign local_bb1_var_[60] = local_bb1_mul[31];
assign local_bb1_var_[61] = local_bb1_mul[31];
assign local_bb1_var_[62] = local_bb1_mul[31];
assign local_bb1_var_[63] = local_bb1_mul[31];
assign local_bb1_var_[31:0] = local_bb1_mul;
assign local_bb1_var__valid_out = local_bb1_var__inputs_ready;
assign local_bb1_var__stall_local = local_bb1_var__stall_in;
assign local_bb1_mul_stall_in = (|local_bb1_var__stall_local);

// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_bb1_var__reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_1_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb1_var__valid_out & rnode_1to4_input_global_id_0_0_valid_out_NO_SHIFT_REG & rnode_1to4_input_global_id_1_0_valid_out_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(stall_in) | ~(branch_node_valid_out_NO_SHIFT_REG));
assign local_bb1_var__stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to4_input_global_id_0_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_1to4_input_global_id_1_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_bb1_var_ = lvb_bb1_var__reg_NO_SHIFT_REG;
assign lvb_input_global_id_0 = lvb_input_global_id_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1 = lvb_input_global_id_1_reg_NO_SHIFT_REG;
assign valid_out = branch_node_valid_out_NO_SHIFT_REG;
assign combined_branch_stall_in_signal = stall_in;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
		lvb_bb1_var__reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_1_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_bb1_var__reg_NO_SHIFT_REG <= local_bb1_var_;
			lvb_input_global_id_0_reg_NO_SHIFT_REG <= rnode_1to4_input_global_id_0_0_NO_SHIFT_REG;
			lvb_input_global_id_1_reg_NO_SHIFT_REG <= rnode_1to4_input_global_id_1_0_NO_SHIFT_REG;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

module Matmul_basic_block_2
	(
		input 		clock,
		input 		resetn,
		input [63:0] 		input_m1r,
		input [63:0] 		input_m1i,
		input [31:0] 		input_col_m2,
		input [31:0] 		input_c1f2,
		input [63:0] 		input_m2r,
		input [63:0] 		input_m2i,
		input 		input_wii_cmp3,
		input 		input_wii_cmp3_NEG,
		input 		valid_in_0,
		output 		stall_out_0,
		input [63:0] 		input_var__0,
		input [63:0] 		input_indvars_iv_0,
		input [31:0] 		input_tmpi_06_0,
		input [31:0] 		input_tmpr_05_0,
		input [31:0] 		input_global_id_0_0,
		input [31:0] 		input_global_id_1_0,
		input 		valid_in_1,
		output 		stall_out_1,
		input [63:0] 		input_var__1,
		input [63:0] 		input_indvars_iv_1,
		input [31:0] 		input_tmpi_06_1,
		input [31:0] 		input_tmpr_05_1,
		input [31:0] 		input_global_id_0_1,
		input [31:0] 		input_global_id_1_1,
		output 		valid_out_0,
		input 		stall_in_0,
		output [63:0] 		lvb_var__0,
		output [63:0] 		lvb_bb2_indvars_iv_next_1_0,
		output 		lvb_bb2_exitcond_0,
		output [159:0] 		lvb_bb2_c0_exit_c0_exi4_0,
		output [31:0] 		lvb_bb2_c0_exe3_0,
		output [31:0] 		lvb_bb2_c0_exe4_0,
		output [31:0] 		lvb_input_global_id_0_0,
		output [31:0] 		lvb_input_global_id_1_0,
		output 		valid_out_1,
		input 		stall_in_1,
		output [63:0] 		lvb_var__1,
		output [63:0] 		lvb_bb2_indvars_iv_next_1_1,
		output 		lvb_bb2_exitcond_1,
		output [159:0] 		lvb_bb2_c0_exit_c0_exi4_1,
		output [31:0] 		lvb_bb2_c0_exe3_1,
		output [31:0] 		lvb_bb2_c0_exe4_1,
		output [31:0] 		lvb_input_global_id_0_1,
		output [31:0] 		lvb_input_global_id_1_1,
		input [31:0] 		workgroup_size,
		input 		start,
		input [255:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_readdata,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_readdatavalid,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_waitrequest,
		output [29:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_address,
		output 		avm_local_bb2_ld_memcoalesce_m1r_load_0_read,
		output 		avm_local_bb2_ld_memcoalesce_m1r_load_0_write,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_writeack,
		output [255:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_writedata,
		output [31:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_byteenable,
		output [4:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_burstcount,
		output 		local_bb2_ld_memcoalesce_m1r_load_0_active,
		input 		clock2x,
		input [255:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_readdata,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_readdatavalid,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_waitrequest,
		output [29:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_address,
		output 		avm_local_bb2_ld_memcoalesce_m1i_load_0_read,
		output 		avm_local_bb2_ld_memcoalesce_m1i_load_0_write,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_writeack,
		output [255:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_writedata,
		output [31:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_byteenable,
		output [4:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_burstcount,
		output 		local_bb2_ld_memcoalesce_m1i_load_0_active,
		input [255:0] 		avm_local_bb2_ld__readdata,
		input 		avm_local_bb2_ld__readdatavalid,
		input 		avm_local_bb2_ld__waitrequest,
		output [29:0] 		avm_local_bb2_ld__address,
		output 		avm_local_bb2_ld__read,
		output 		avm_local_bb2_ld__write,
		input 		avm_local_bb2_ld__writeack,
		output [255:0] 		avm_local_bb2_ld__writedata,
		output [31:0] 		avm_local_bb2_ld__byteenable,
		output [4:0] 		avm_local_bb2_ld__burstcount,
		output 		local_bb2_ld__active,
		input [255:0] 		avm_local_bb2_ld__u1_readdata,
		input 		avm_local_bb2_ld__u1_readdatavalid,
		input 		avm_local_bb2_ld__u1_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u1_address,
		output 		avm_local_bb2_ld__u1_read,
		output 		avm_local_bb2_ld__u1_write,
		input 		avm_local_bb2_ld__u1_writeack,
		output [255:0] 		avm_local_bb2_ld__u1_writedata,
		output [31:0] 		avm_local_bb2_ld__u1_byteenable,
		output [4:0] 		avm_local_bb2_ld__u1_burstcount,
		output 		local_bb2_ld__u1_active,
		input [255:0] 		avm_local_bb2_ld__u2_readdata,
		input 		avm_local_bb2_ld__u2_readdatavalid,
		input 		avm_local_bb2_ld__u2_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u2_address,
		output 		avm_local_bb2_ld__u2_read,
		output 		avm_local_bb2_ld__u2_write,
		input 		avm_local_bb2_ld__u2_writeack,
		output [255:0] 		avm_local_bb2_ld__u2_writedata,
		output [31:0] 		avm_local_bb2_ld__u2_byteenable,
		output [4:0] 		avm_local_bb2_ld__u2_burstcount,
		output 		local_bb2_ld__u2_active,
		input [255:0] 		avm_local_bb2_ld__u3_readdata,
		input 		avm_local_bb2_ld__u3_readdatavalid,
		input 		avm_local_bb2_ld__u3_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u3_address,
		output 		avm_local_bb2_ld__u3_read,
		output 		avm_local_bb2_ld__u3_write,
		input 		avm_local_bb2_ld__u3_writeack,
		output [255:0] 		avm_local_bb2_ld__u3_writedata,
		output [31:0] 		avm_local_bb2_ld__u3_byteenable,
		output [4:0] 		avm_local_bb2_ld__u3_burstcount,
		output 		local_bb2_ld__u3_active
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((valid_in_0 & valid_in_1) & ~((stall_out_0 | stall_out_1)));
assign _exit = ((valid_out_0 & valid_out_1) & ~((stall_in_0 | stall_in_1)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_node_stall_in_6;
 reg merge_node_valid_out_6_NO_SHIFT_REG;
wire merge_node_stall_in_7;
 reg merge_node_valid_out_7_NO_SHIFT_REG;
wire merge_node_stall_in_8;
 reg merge_node_valid_out_8_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_var__0_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_tmpi_06_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_tmpr_05_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_0_staging_reg_NO_SHIFT_REG;
 reg [63:0] local_lvm_var__NO_SHIFT_REG;
 reg [63:0] local_lvm_indvars_iv_NO_SHIFT_REG;
 reg [31:0] local_lvm_tmpi_06_NO_SHIFT_REG;
 reg [31:0] local_lvm_tmpr_05_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_var__1_staging_reg_NO_SHIFT_REG;
 reg [63:0] input_indvars_iv_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_tmpi_06_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_tmpr_05_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_1_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_1_staging_reg_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG) | (merge_node_stall_in_6 & merge_node_valid_out_6_NO_SHIFT_REG) | (merge_node_stall_in_7 & merge_node_valid_out_7_NO_SHIFT_REG) | (merge_node_stall_in_8 & merge_node_valid_out_8_NO_SHIFT_REG));
assign stall_out_0 = merge_node_valid_in_0_staging_reg_NO_SHIFT_REG;
assign stall_out_1 = merge_node_valid_in_1_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_0_staging_reg_NO_SHIFT_REG | valid_in_0))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		if ((merge_node_valid_in_1_staging_reg_NO_SHIFT_REG | valid_in_1))
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b1;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
		end
		else
		begin
			merge_block_selector_NO_SHIFT_REG = 1'b0;
			is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_var__0_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_tmpi_06_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_tmpr_05_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_0_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_0_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		input_var__1_staging_reg_NO_SHIFT_REG <= 'x;
		input_indvars_iv_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_tmpi_06_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_tmpr_05_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_0_1_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_0_staging_reg_NO_SHIFT_REG))
			begin
				input_var__0_staging_reg_NO_SHIFT_REG <= input_var__0;
				input_indvars_iv_0_staging_reg_NO_SHIFT_REG <= input_indvars_iv_0;
				input_tmpi_06_0_staging_reg_NO_SHIFT_REG <= input_tmpi_06_0;
				input_tmpr_05_0_staging_reg_NO_SHIFT_REG <= input_tmpr_05_0;
				input_global_id_0_0_staging_reg_NO_SHIFT_REG <= input_global_id_0_0;
				input_global_id_1_0_staging_reg_NO_SHIFT_REG <= input_global_id_1_0;
				merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= valid_in_0;
			end
		end
		else
		begin
			merge_node_valid_in_0_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
		if (((merge_block_selector_NO_SHIFT_REG != 1'b1) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_1_staging_reg_NO_SHIFT_REG))
			begin
				input_var__1_staging_reg_NO_SHIFT_REG <= input_var__1;
				input_indvars_iv_1_staging_reg_NO_SHIFT_REG <= input_indvars_iv_1;
				input_tmpi_06_1_staging_reg_NO_SHIFT_REG <= input_tmpi_06_1;
				input_tmpr_05_1_staging_reg_NO_SHIFT_REG <= input_tmpr_05_1;
				input_global_id_0_1_staging_reg_NO_SHIFT_REG <= input_global_id_0_1;
				input_global_id_1_1_staging_reg_NO_SHIFT_REG <= input_global_id_1_1;
				merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= valid_in_1;
			end
		end
		else
		begin
			merge_node_valid_in_1_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_0_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_var__NO_SHIFT_REG <= input_var__0_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv_NO_SHIFT_REG <= input_indvars_iv_0_staging_reg_NO_SHIFT_REG;
					local_lvm_tmpi_06_NO_SHIFT_REG <= input_tmpi_06_0_staging_reg_NO_SHIFT_REG;
					local_lvm_tmpr_05_NO_SHIFT_REG <= input_tmpr_05_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_0_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_var__NO_SHIFT_REG <= input_var__0;
					local_lvm_indvars_iv_NO_SHIFT_REG <= input_indvars_iv_0;
					local_lvm_tmpi_06_NO_SHIFT_REG <= input_tmpi_06_0;
					local_lvm_tmpr_05_NO_SHIFT_REG <= input_tmpr_05_0;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_0;
				end
			end

			1'b1:
			begin
				if (merge_node_valid_in_1_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_var__NO_SHIFT_REG <= input_var__1_staging_reg_NO_SHIFT_REG;
					local_lvm_indvars_iv_NO_SHIFT_REG <= input_indvars_iv_1_staging_reg_NO_SHIFT_REG;
					local_lvm_tmpi_06_NO_SHIFT_REG <= input_tmpi_06_1_staging_reg_NO_SHIFT_REG;
					local_lvm_tmpr_05_NO_SHIFT_REG <= input_tmpr_05_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_1_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_var__NO_SHIFT_REG <= input_var__1;
					local_lvm_indvars_iv_NO_SHIFT_REG <= input_indvars_iv_1;
					local_lvm_tmpi_06_NO_SHIFT_REG <= input_tmpi_06_1;
					local_lvm_tmpr_05_NO_SHIFT_REG <= input_tmpr_05_1;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_1;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_6_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_7_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_8_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_6))
			begin
				merge_node_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_7))
			begin
				merge_node_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_8))
			begin
				merge_node_valid_out_8_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_indvars_iv_next10_stall_local;
wire [63:0] local_bb2_indvars_iv_next10;

assign local_bb2_indvars_iv_next10 = (local_lvm_indvars_iv_NO_SHIFT_REG | 64'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__valid_out;
wire local_bb2_var__stall_in;
wire local_bb2_var__inputs_ready;
wire local_bb2_var__stall_local;
wire [31:0] local_bb2_var_;

assign local_bb2_var__inputs_ready = merge_node_valid_out_1_NO_SHIFT_REG;
assign local_bb2_var_ = local_lvm_indvars_iv_NO_SHIFT_REG[31:0];
assign local_bb2_var__valid_out = local_bb2_var__inputs_ready;
assign local_bb2_var__stall_local = local_bb2_var__stall_in;
assign merge_node_stall_in_1 = (|local_bb2_var__stall_local);

// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_1to5_cmp3_NEG_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_stall_in_3_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_valid_out_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_stall_in_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_cmp3_NEG_0_stall_out_reg_5_NO_SHIFT_REG;

acl_multi_fanout_adaptor rnode_1to5_cmp3_NEG_0_reg_5_fanout_adaptor (
	.clock(clock),
	.resetn(resetn),
	.data_in(),
	.valid_in(rnode_1to5_cmp3_NEG_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_1to5_cmp3_NEG_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.data_out(),
	.valid_out({rnode_1to5_cmp3_NEG_0_valid_out_0_NO_SHIFT_REG, rnode_1to5_cmp3_NEG_0_valid_out_1_NO_SHIFT_REG, rnode_1to5_cmp3_NEG_0_valid_out_2_NO_SHIFT_REG, rnode_1to5_cmp3_NEG_0_valid_out_3_NO_SHIFT_REG}),
	.stall_in({rnode_1to5_cmp3_NEG_0_stall_in_0_NO_SHIFT_REG, rnode_1to5_cmp3_NEG_0_stall_in_1_NO_SHIFT_REG, rnode_1to5_cmp3_NEG_0_stall_in_2_NO_SHIFT_REG, rnode_1to5_cmp3_NEG_0_stall_in_3_NO_SHIFT_REG})
);

defparam rnode_1to5_cmp3_NEG_0_reg_5_fanout_adaptor.DATA_WIDTH = 0;
defparam rnode_1to5_cmp3_NEG_0_reg_5_fanout_adaptor.NUM_FANOUTS = 4;

acl_data_fifo rnode_1to5_cmp3_NEG_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to5_cmp3_NEG_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to5_cmp3_NEG_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_1to5_cmp3_NEG_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_1to5_cmp3_NEG_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(),
	.data_out()
);

defparam rnode_1to5_cmp3_NEG_0_reg_5_fifo.DEPTH = 5;
defparam rnode_1to5_cmp3_NEG_0_reg_5_fifo.DATA_WIDTH = 0;
defparam rnode_1to5_cmp3_NEG_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to5_cmp3_NEG_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_1to5_cmp3_NEG_0_reg_5_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_2_NO_SHIFT_REG;
assign merge_node_stall_in_2 = rnode_1to5_cmp3_NEG_0_stall_out_reg_5_NO_SHIFT_REG;

// Register node:
//  * latency = 163
//  * capacity = 163
 logic rnode_1to164_tmpr_05_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to164_tmpr_05_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to164_tmpr_05_0_NO_SHIFT_REG;
 logic rnode_1to164_tmpr_05_0_reg_164_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to164_tmpr_05_0_reg_164_NO_SHIFT_REG;
 logic rnode_1to164_tmpr_05_0_valid_out_reg_164_NO_SHIFT_REG;
 logic rnode_1to164_tmpr_05_0_stall_in_reg_164_NO_SHIFT_REG;
 logic rnode_1to164_tmpr_05_0_stall_out_reg_164_NO_SHIFT_REG;

acl_data_fifo rnode_1to164_tmpr_05_0_reg_164_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to164_tmpr_05_0_reg_164_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to164_tmpr_05_0_stall_in_reg_164_NO_SHIFT_REG),
	.valid_out(rnode_1to164_tmpr_05_0_valid_out_reg_164_NO_SHIFT_REG),
	.stall_out(rnode_1to164_tmpr_05_0_stall_out_reg_164_NO_SHIFT_REG),
	.data_in(local_lvm_tmpr_05_NO_SHIFT_REG),
	.data_out(rnode_1to164_tmpr_05_0_reg_164_NO_SHIFT_REG)
);

defparam rnode_1to164_tmpr_05_0_reg_164_fifo.DEPTH = 164;
defparam rnode_1to164_tmpr_05_0_reg_164_fifo.DATA_WIDTH = 32;
defparam rnode_1to164_tmpr_05_0_reg_164_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to164_tmpr_05_0_reg_164_fifo.IMPL = "ram";

assign rnode_1to164_tmpr_05_0_reg_164_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_3_NO_SHIFT_REG;
assign merge_node_stall_in_3 = rnode_1to164_tmpr_05_0_stall_out_reg_164_NO_SHIFT_REG;
assign rnode_1to164_tmpr_05_0_NO_SHIFT_REG = rnode_1to164_tmpr_05_0_reg_164_NO_SHIFT_REG;
assign rnode_1to164_tmpr_05_0_stall_in_reg_164_NO_SHIFT_REG = rnode_1to164_tmpr_05_0_stall_in_NO_SHIFT_REG;
assign rnode_1to164_tmpr_05_0_valid_out_NO_SHIFT_REG = rnode_1to164_tmpr_05_0_valid_out_reg_164_NO_SHIFT_REG;

// Register node:
//  * latency = 163
//  * capacity = 163
 logic rnode_1to164_tmpi_06_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to164_tmpi_06_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to164_tmpi_06_0_NO_SHIFT_REG;
 logic rnode_1to164_tmpi_06_0_reg_164_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to164_tmpi_06_0_reg_164_NO_SHIFT_REG;
 logic rnode_1to164_tmpi_06_0_valid_out_reg_164_NO_SHIFT_REG;
 logic rnode_1to164_tmpi_06_0_stall_in_reg_164_NO_SHIFT_REG;
 logic rnode_1to164_tmpi_06_0_stall_out_reg_164_NO_SHIFT_REG;

acl_data_fifo rnode_1to164_tmpi_06_0_reg_164_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to164_tmpi_06_0_reg_164_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to164_tmpi_06_0_stall_in_reg_164_NO_SHIFT_REG),
	.valid_out(rnode_1to164_tmpi_06_0_valid_out_reg_164_NO_SHIFT_REG),
	.stall_out(rnode_1to164_tmpi_06_0_stall_out_reg_164_NO_SHIFT_REG),
	.data_in(local_lvm_tmpi_06_NO_SHIFT_REG),
	.data_out(rnode_1to164_tmpi_06_0_reg_164_NO_SHIFT_REG)
);

defparam rnode_1to164_tmpi_06_0_reg_164_fifo.DEPTH = 164;
defparam rnode_1to164_tmpi_06_0_reg_164_fifo.DATA_WIDTH = 32;
defparam rnode_1to164_tmpi_06_0_reg_164_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to164_tmpi_06_0_reg_164_fifo.IMPL = "ram";

assign rnode_1to164_tmpi_06_0_reg_164_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_4_NO_SHIFT_REG;
assign merge_node_stall_in_4 = rnode_1to164_tmpi_06_0_stall_out_reg_164_NO_SHIFT_REG;
assign rnode_1to164_tmpi_06_0_NO_SHIFT_REG = rnode_1to164_tmpi_06_0_reg_164_NO_SHIFT_REG;
assign rnode_1to164_tmpi_06_0_stall_in_reg_164_NO_SHIFT_REG = rnode_1to164_tmpi_06_0_stall_in_NO_SHIFT_REG;
assign rnode_1to164_tmpi_06_0_valid_out_NO_SHIFT_REG = rnode_1to164_tmpi_06_0_valid_out_reg_164_NO_SHIFT_REG;

// Register node:
//  * latency = 194
//  * capacity = 194
 logic rnode_1to195_input_global_id_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to195_input_global_id_1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to195_input_global_id_1_0_NO_SHIFT_REG;
 logic rnode_1to195_input_global_id_1_0_reg_195_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to195_input_global_id_1_0_reg_195_NO_SHIFT_REG;
 logic rnode_1to195_input_global_id_1_0_valid_out_reg_195_NO_SHIFT_REG;
 logic rnode_1to195_input_global_id_1_0_stall_in_reg_195_NO_SHIFT_REG;
 logic rnode_1to195_input_global_id_1_0_stall_out_reg_195_NO_SHIFT_REG;

acl_data_fifo rnode_1to195_input_global_id_1_0_reg_195_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to195_input_global_id_1_0_reg_195_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to195_input_global_id_1_0_stall_in_reg_195_NO_SHIFT_REG),
	.valid_out(rnode_1to195_input_global_id_1_0_valid_out_reg_195_NO_SHIFT_REG),
	.stall_out(rnode_1to195_input_global_id_1_0_stall_out_reg_195_NO_SHIFT_REG),
	.data_in(local_lvm_input_global_id_1_NO_SHIFT_REG),
	.data_out(rnode_1to195_input_global_id_1_0_reg_195_NO_SHIFT_REG)
);

defparam rnode_1to195_input_global_id_1_0_reg_195_fifo.DEPTH = 195;
defparam rnode_1to195_input_global_id_1_0_reg_195_fifo.DATA_WIDTH = 32;
defparam rnode_1to195_input_global_id_1_0_reg_195_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to195_input_global_id_1_0_reg_195_fifo.IMPL = "ram";

assign rnode_1to195_input_global_id_1_0_reg_195_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_5_NO_SHIFT_REG;
assign merge_node_stall_in_5 = rnode_1to195_input_global_id_1_0_stall_out_reg_195_NO_SHIFT_REG;
assign rnode_1to195_input_global_id_1_0_NO_SHIFT_REG = rnode_1to195_input_global_id_1_0_reg_195_NO_SHIFT_REG;
assign rnode_1to195_input_global_id_1_0_stall_in_reg_195_NO_SHIFT_REG = rnode_1to195_input_global_id_1_0_stall_in_NO_SHIFT_REG;
assign rnode_1to195_input_global_id_1_0_valid_out_NO_SHIFT_REG = rnode_1to195_input_global_id_1_0_valid_out_reg_195_NO_SHIFT_REG;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_indvars_iv_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to4_indvars_iv_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_1to4_indvars_iv_0_NO_SHIFT_REG;
 logic rnode_1to4_indvars_iv_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to4_indvars_iv_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_1to4_indvars_iv_1_NO_SHIFT_REG;
 logic rnode_1to4_indvars_iv_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to4_indvars_iv_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_indvars_iv_0_valid_out_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_indvars_iv_0_stall_in_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_indvars_iv_0_stall_out_reg_4_NO_SHIFT_REG;
 logic [63:0] rnode_1to4_indvars_iv_0_reg_4_NO_SHIFT_REG_fa;

acl_multi_fanout_adaptor rnode_1to4_indvars_iv_0_reg_4_fanout_adaptor (
	.clock(clock),
	.resetn(resetn),
	.data_in(rnode_1to4_indvars_iv_0_reg_4_NO_SHIFT_REG),
	.valid_in(rnode_1to4_indvars_iv_0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_indvars_iv_0_stall_in_0_reg_4_NO_SHIFT_REG),
	.data_out(rnode_1to4_indvars_iv_0_reg_4_NO_SHIFT_REG_fa),
	.valid_out({rnode_1to4_indvars_iv_0_valid_out_0_NO_SHIFT_REG, rnode_1to4_indvars_iv_0_valid_out_1_NO_SHIFT_REG}),
	.stall_in({rnode_1to4_indvars_iv_0_stall_in_0_NO_SHIFT_REG, rnode_1to4_indvars_iv_0_stall_in_1_NO_SHIFT_REG})
);

defparam rnode_1to4_indvars_iv_0_reg_4_fanout_adaptor.DATA_WIDTH = 64;
defparam rnode_1to4_indvars_iv_0_reg_4_fanout_adaptor.NUM_FANOUTS = 2;

acl_data_fifo rnode_1to4_indvars_iv_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_indvars_iv_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_indvars_iv_0_stall_in_0_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_indvars_iv_0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_indvars_iv_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_lvm_indvars_iv_NO_SHIFT_REG),
	.data_out(rnode_1to4_indvars_iv_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_indvars_iv_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_indvars_iv_0_reg_4_fifo.DATA_WIDTH = 64;
defparam rnode_1to4_indvars_iv_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_indvars_iv_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_indvars_iv_0_reg_4_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_6_NO_SHIFT_REG;
assign merge_node_stall_in_6 = rnode_1to4_indvars_iv_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_indvars_iv_0_NO_SHIFT_REG = rnode_1to4_indvars_iv_0_reg_4_NO_SHIFT_REG_fa;
assign rnode_1to4_indvars_iv_1_NO_SHIFT_REG = rnode_1to4_indvars_iv_0_reg_4_NO_SHIFT_REG_fa;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_var__0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to4_var__0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_1to4_var__0_NO_SHIFT_REG;
 logic rnode_1to4_var__0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to4_var__0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_1to4_var__1_NO_SHIFT_REG;
 logic rnode_1to4_var__0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_1to4_var__0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_var__0_valid_out_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_var__0_stall_in_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_var__0_stall_out_reg_4_NO_SHIFT_REG;
 logic [63:0] rnode_1to4_var__0_reg_4_NO_SHIFT_REG_fa;

acl_multi_fanout_adaptor rnode_1to4_var__0_reg_4_fanout_adaptor (
	.clock(clock),
	.resetn(resetn),
	.data_in(rnode_1to4_var__0_reg_4_NO_SHIFT_REG),
	.valid_in(rnode_1to4_var__0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_var__0_stall_in_0_reg_4_NO_SHIFT_REG),
	.data_out(rnode_1to4_var__0_reg_4_NO_SHIFT_REG_fa),
	.valid_out({rnode_1to4_var__0_valid_out_0_NO_SHIFT_REG, rnode_1to4_var__0_valid_out_1_NO_SHIFT_REG}),
	.stall_in({rnode_1to4_var__0_stall_in_0_NO_SHIFT_REG, rnode_1to4_var__0_stall_in_1_NO_SHIFT_REG})
);

defparam rnode_1to4_var__0_reg_4_fanout_adaptor.DATA_WIDTH = 64;
defparam rnode_1to4_var__0_reg_4_fanout_adaptor.NUM_FANOUTS = 2;

acl_data_fifo rnode_1to4_var__0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_var__0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_var__0_stall_in_0_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_var__0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_var__0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_lvm_var__NO_SHIFT_REG),
	.data_out(rnode_1to4_var__0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_var__0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_var__0_reg_4_fifo.DATA_WIDTH = 64;
defparam rnode_1to4_var__0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_var__0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_var__0_reg_4_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_7_NO_SHIFT_REG;
assign merge_node_stall_in_7 = rnode_1to4_var__0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_var__0_NO_SHIFT_REG = rnode_1to4_var__0_reg_4_NO_SHIFT_REG_fa;
assign rnode_1to4_var__1_NO_SHIFT_REG = rnode_1to4_var__0_reg_4_NO_SHIFT_REG_fa;

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_input_global_id_0_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_1_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_2_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG_fa;

acl_multi_fanout_adaptor rnode_1to4_input_global_id_0_0_reg_4_fanout_adaptor (
	.clock(clock),
	.resetn(resetn),
	.data_in(rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG),
	.valid_in(rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_input_global_id_0_0_stall_in_0_reg_4_NO_SHIFT_REG),
	.data_out(rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG_fa),
	.valid_out({rnode_1to4_input_global_id_0_0_valid_out_0_NO_SHIFT_REG, rnode_1to4_input_global_id_0_0_valid_out_1_NO_SHIFT_REG, rnode_1to4_input_global_id_0_0_valid_out_2_NO_SHIFT_REG}),
	.stall_in({rnode_1to4_input_global_id_0_0_stall_in_0_NO_SHIFT_REG, rnode_1to4_input_global_id_0_0_stall_in_1_NO_SHIFT_REG, rnode_1to4_input_global_id_0_0_stall_in_2_NO_SHIFT_REG})
);

defparam rnode_1to4_input_global_id_0_0_reg_4_fanout_adaptor.DATA_WIDTH = 32;
defparam rnode_1to4_input_global_id_0_0_reg_4_fanout_adaptor.NUM_FANOUTS = 3;

acl_data_fifo rnode_1to4_input_global_id_0_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_input_global_id_0_0_stall_in_0_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_input_global_id_0_0_valid_out_0_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_lvm_input_global_id_0_NO_SHIFT_REG),
	.data_out(rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_8_NO_SHIFT_REG;
assign merge_node_stall_in_8 = rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG_fa;
assign rnode_1to4_input_global_id_0_1_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG_fa;
assign rnode_1to4_input_global_id_0_2_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG_fa;

// This section implements an unregistered operation.
// 
wire local_bb2_lftr_wideiv_stall_local;
wire [31:0] local_bb2_lftr_wideiv;

assign local_bb2_lftr_wideiv = local_bb2_indvars_iv_next10[31:0];

// This section implements a registered operation.
// 
wire local_bb2_mul4_inputs_ready;
 reg local_bb2_mul4_valid_out_NO_SHIFT_REG;
wire local_bb2_mul4_stall_in;
wire local_bb2_mul4_output_regs_ready;
wire [31:0] local_bb2_mul4;
 reg local_bb2_mul4_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul4_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul4_causedstall;

acl_int_mult32s_s5 int_module_local_bb2_mul4 (
	.clock(clock),
	.dataa(local_bb2_var_),
	.datab(input_col_m2),
	.enable(local_bb2_mul4_output_regs_ready),
	.result(local_bb2_mul4)
);

defparam int_module_local_bb2_mul4.INPUT1_WIDTH = 32;
defparam int_module_local_bb2_mul4.INPUT2_WIDTH = 32;

assign local_bb2_mul4_inputs_ready = local_bb2_var__valid_out;
assign local_bb2_mul4_output_regs_ready = (&(~(local_bb2_mul4_valid_out_NO_SHIFT_REG) | ~(local_bb2_mul4_stall_in)));
assign local_bb2_var__stall_in = (~(local_bb2_mul4_output_regs_ready) | ~(local_bb2_mul4_inputs_ready));
assign local_bb2_mul4_causedstall = (local_bb2_mul4_inputs_ready && (~(local_bb2_mul4_output_regs_ready) && !(~(local_bb2_mul4_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul4_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul4_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul4_output_regs_ready)
		begin
			local_bb2_mul4_valid_pipe_0_NO_SHIFT_REG <= local_bb2_mul4_inputs_ready;
			local_bb2_mul4_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul4_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul4_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul4_output_regs_ready)
		begin
			local_bb2_mul4_valid_out_NO_SHIFT_REG <= local_bb2_mul4_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb2_mul4_stall_in))
			begin
				local_bb2_mul4_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_164to165_tmpr_05_0_valid_out_NO_SHIFT_REG;
 logic rnode_164to165_tmpr_05_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_164to165_tmpr_05_0_NO_SHIFT_REG;
 logic rnode_164to165_tmpr_05_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_164to165_tmpr_05_0_reg_165_NO_SHIFT_REG;
 logic rnode_164to165_tmpr_05_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_164to165_tmpr_05_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_164to165_tmpr_05_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_164to165_tmpr_05_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_164to165_tmpr_05_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_164to165_tmpr_05_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_164to165_tmpr_05_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_164to165_tmpr_05_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(rnode_1to164_tmpr_05_0_NO_SHIFT_REG),
	.data_out(rnode_164to165_tmpr_05_0_reg_165_NO_SHIFT_REG)
);

defparam rnode_164to165_tmpr_05_0_reg_165_fifo.DEPTH = 2;
defparam rnode_164to165_tmpr_05_0_reg_165_fifo.DATA_WIDTH = 32;
defparam rnode_164to165_tmpr_05_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_164to165_tmpr_05_0_reg_165_fifo.IMPL = "ll_reg";

assign rnode_164to165_tmpr_05_0_reg_165_inputs_ready_NO_SHIFT_REG = rnode_1to164_tmpr_05_0_valid_out_NO_SHIFT_REG;
assign rnode_1to164_tmpr_05_0_stall_in_NO_SHIFT_REG = rnode_164to165_tmpr_05_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_164to165_tmpr_05_0_NO_SHIFT_REG = rnode_164to165_tmpr_05_0_reg_165_NO_SHIFT_REG;
assign rnode_164to165_tmpr_05_0_stall_in_reg_165_NO_SHIFT_REG = rnode_164to165_tmpr_05_0_stall_in_NO_SHIFT_REG;
assign rnode_164to165_tmpr_05_0_valid_out_NO_SHIFT_REG = rnode_164to165_tmpr_05_0_valid_out_reg_165_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_164to165_tmpi_06_0_valid_out_NO_SHIFT_REG;
 logic rnode_164to165_tmpi_06_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_164to165_tmpi_06_0_NO_SHIFT_REG;
 logic rnode_164to165_tmpi_06_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_164to165_tmpi_06_0_reg_165_NO_SHIFT_REG;
 logic rnode_164to165_tmpi_06_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_164to165_tmpi_06_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_164to165_tmpi_06_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_164to165_tmpi_06_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_164to165_tmpi_06_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_164to165_tmpi_06_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_164to165_tmpi_06_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_164to165_tmpi_06_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(rnode_1to164_tmpi_06_0_NO_SHIFT_REG),
	.data_out(rnode_164to165_tmpi_06_0_reg_165_NO_SHIFT_REG)
);

defparam rnode_164to165_tmpi_06_0_reg_165_fifo.DEPTH = 2;
defparam rnode_164to165_tmpi_06_0_reg_165_fifo.DATA_WIDTH = 32;
defparam rnode_164to165_tmpi_06_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_164to165_tmpi_06_0_reg_165_fifo.IMPL = "ll_reg";

assign rnode_164to165_tmpi_06_0_reg_165_inputs_ready_NO_SHIFT_REG = rnode_1to164_tmpi_06_0_valid_out_NO_SHIFT_REG;
assign rnode_1to164_tmpi_06_0_stall_in_NO_SHIFT_REG = rnode_164to165_tmpi_06_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_164to165_tmpi_06_0_NO_SHIFT_REG = rnode_164to165_tmpi_06_0_reg_165_NO_SHIFT_REG;
assign rnode_164to165_tmpi_06_0_stall_in_reg_165_NO_SHIFT_REG = rnode_164to165_tmpi_06_0_stall_in_NO_SHIFT_REG;
assign rnode_164to165_tmpi_06_0_valid_out_NO_SHIFT_REG = rnode_164to165_tmpi_06_0_valid_out_reg_165_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_195to196_input_global_id_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_195to196_input_global_id_1_0_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_1_0_reg_196_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_195to196_input_global_id_1_0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_1_0_valid_out_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_1_0_stall_in_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_1_0_stall_out_reg_196_NO_SHIFT_REG;

acl_data_fifo rnode_195to196_input_global_id_1_0_reg_196_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_195to196_input_global_id_1_0_reg_196_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_195to196_input_global_id_1_0_stall_in_reg_196_NO_SHIFT_REG),
	.valid_out(rnode_195to196_input_global_id_1_0_valid_out_reg_196_NO_SHIFT_REG),
	.stall_out(rnode_195to196_input_global_id_1_0_stall_out_reg_196_NO_SHIFT_REG),
	.data_in(rnode_1to195_input_global_id_1_0_NO_SHIFT_REG),
	.data_out(rnode_195to196_input_global_id_1_0_reg_196_NO_SHIFT_REG)
);

defparam rnode_195to196_input_global_id_1_0_reg_196_fifo.DEPTH = 2;
defparam rnode_195to196_input_global_id_1_0_reg_196_fifo.DATA_WIDTH = 32;
defparam rnode_195to196_input_global_id_1_0_reg_196_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_195to196_input_global_id_1_0_reg_196_fifo.IMPL = "ll_reg";

assign rnode_195to196_input_global_id_1_0_reg_196_inputs_ready_NO_SHIFT_REG = rnode_1to195_input_global_id_1_0_valid_out_NO_SHIFT_REG;
assign rnode_1to195_input_global_id_1_0_stall_in_NO_SHIFT_REG = rnode_195to196_input_global_id_1_0_stall_out_reg_196_NO_SHIFT_REG;
assign rnode_195to196_input_global_id_1_0_NO_SHIFT_REG = rnode_195to196_input_global_id_1_0_reg_196_NO_SHIFT_REG;
assign rnode_195to196_input_global_id_1_0_stall_in_reg_196_NO_SHIFT_REG = rnode_195to196_input_global_id_1_0_stall_in_NO_SHIFT_REG;
assign rnode_195to196_input_global_id_1_0_valid_out_NO_SHIFT_REG = rnode_195to196_input_global_id_1_0_valid_out_reg_196_NO_SHIFT_REG;

// Register node:
//  * latency = 190
//  * capacity = 190
 logic rnode_4to194_indvars_iv_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to194_indvars_iv_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_4to194_indvars_iv_0_NO_SHIFT_REG;
 logic rnode_4to194_indvars_iv_0_reg_194_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_4to194_indvars_iv_0_reg_194_NO_SHIFT_REG;
 logic rnode_4to194_indvars_iv_0_valid_out_reg_194_NO_SHIFT_REG;
 logic rnode_4to194_indvars_iv_0_stall_in_reg_194_NO_SHIFT_REG;
 logic rnode_4to194_indvars_iv_0_stall_out_reg_194_NO_SHIFT_REG;

acl_data_fifo rnode_4to194_indvars_iv_0_reg_194_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to194_indvars_iv_0_reg_194_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to194_indvars_iv_0_stall_in_reg_194_NO_SHIFT_REG),
	.valid_out(rnode_4to194_indvars_iv_0_valid_out_reg_194_NO_SHIFT_REG),
	.stall_out(rnode_4to194_indvars_iv_0_stall_out_reg_194_NO_SHIFT_REG),
	.data_in(rnode_1to4_indvars_iv_1_NO_SHIFT_REG),
	.data_out(rnode_4to194_indvars_iv_0_reg_194_NO_SHIFT_REG)
);

defparam rnode_4to194_indvars_iv_0_reg_194_fifo.DEPTH = 191;
defparam rnode_4to194_indvars_iv_0_reg_194_fifo.DATA_WIDTH = 64;
defparam rnode_4to194_indvars_iv_0_reg_194_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to194_indvars_iv_0_reg_194_fifo.IMPL = "ram";

assign rnode_4to194_indvars_iv_0_reg_194_inputs_ready_NO_SHIFT_REG = rnode_1to4_indvars_iv_0_valid_out_1_NO_SHIFT_REG;
assign rnode_1to4_indvars_iv_0_stall_in_1_NO_SHIFT_REG = rnode_4to194_indvars_iv_0_stall_out_reg_194_NO_SHIFT_REG;
assign rnode_4to194_indvars_iv_0_NO_SHIFT_REG = rnode_4to194_indvars_iv_0_reg_194_NO_SHIFT_REG;
assign rnode_4to194_indvars_iv_0_stall_in_reg_194_NO_SHIFT_REG = rnode_4to194_indvars_iv_0_stall_in_NO_SHIFT_REG;
assign rnode_4to194_indvars_iv_0_valid_out_NO_SHIFT_REG = rnode_4to194_indvars_iv_0_valid_out_reg_194_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u0_valid_out;
wire local_bb2_var__u0_stall_in;
wire local_bb2_var__u0_inputs_ready;
wire local_bb2_var__u0_stall_local;
wire [63:0] local_bb2_var__u0;

assign local_bb2_var__u0_inputs_ready = (rnode_1to4_indvars_iv_0_valid_out_0_NO_SHIFT_REG & rnode_1to4_var__0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_var__u0 = (rnode_1to4_indvars_iv_0_NO_SHIFT_REG + rnode_1to4_var__0_NO_SHIFT_REG);
assign local_bb2_var__u0_valid_out = local_bb2_var__u0_inputs_ready;
assign local_bb2_var__u0_stall_local = local_bb2_var__u0_stall_in;
assign rnode_1to4_indvars_iv_0_stall_in_0_NO_SHIFT_REG = (local_bb2_var__u0_stall_local | ~(local_bb2_var__u0_inputs_ready));
assign rnode_1to4_var__0_stall_in_0_NO_SHIFT_REG = (local_bb2_var__u0_stall_local | ~(local_bb2_var__u0_inputs_ready));

// Register node:
//  * latency = 191
//  * capacity = 191
 logic rnode_4to195_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_4to195_var__0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_4to195_var__0_NO_SHIFT_REG;
 logic rnode_4to195_var__0_reg_195_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_4to195_var__0_reg_195_NO_SHIFT_REG;
 logic rnode_4to195_var__0_valid_out_reg_195_NO_SHIFT_REG;
 logic rnode_4to195_var__0_stall_in_reg_195_NO_SHIFT_REG;
 logic rnode_4to195_var__0_stall_out_reg_195_NO_SHIFT_REG;

acl_data_fifo rnode_4to195_var__0_reg_195_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to195_var__0_reg_195_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to195_var__0_stall_in_reg_195_NO_SHIFT_REG),
	.valid_out(rnode_4to195_var__0_valid_out_reg_195_NO_SHIFT_REG),
	.stall_out(rnode_4to195_var__0_stall_out_reg_195_NO_SHIFT_REG),
	.data_in(rnode_1to4_var__1_NO_SHIFT_REG),
	.data_out(rnode_4to195_var__0_reg_195_NO_SHIFT_REG)
);

defparam rnode_4to195_var__0_reg_195_fifo.DEPTH = 192;
defparam rnode_4to195_var__0_reg_195_fifo.DATA_WIDTH = 64;
defparam rnode_4to195_var__0_reg_195_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to195_var__0_reg_195_fifo.IMPL = "ram";

assign rnode_4to195_var__0_reg_195_inputs_ready_NO_SHIFT_REG = rnode_1to4_var__0_valid_out_1_NO_SHIFT_REG;
assign rnode_1to4_var__0_stall_in_1_NO_SHIFT_REG = rnode_4to195_var__0_stall_out_reg_195_NO_SHIFT_REG;
assign rnode_4to195_var__0_NO_SHIFT_REG = rnode_4to195_var__0_reg_195_NO_SHIFT_REG;
assign rnode_4to195_var__0_stall_in_reg_195_NO_SHIFT_REG = rnode_4to195_var__0_stall_in_NO_SHIFT_REG;
assign rnode_4to195_var__0_valid_out_NO_SHIFT_REG = rnode_4to195_var__0_valid_out_reg_195_NO_SHIFT_REG;

// Register node:
//  * latency = 191
//  * capacity = 191
 logic rnode_4to195_input_global_id_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to195_input_global_id_0_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to195_input_global_id_0_0_NO_SHIFT_REG;
 logic rnode_4to195_input_global_id_0_0_reg_195_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to195_input_global_id_0_0_reg_195_NO_SHIFT_REG;
 logic rnode_4to195_input_global_id_0_0_valid_out_reg_195_NO_SHIFT_REG;
 logic rnode_4to195_input_global_id_0_0_stall_in_reg_195_NO_SHIFT_REG;
 logic rnode_4to195_input_global_id_0_0_stall_out_reg_195_NO_SHIFT_REG;

acl_data_fifo rnode_4to195_input_global_id_0_0_reg_195_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to195_input_global_id_0_0_reg_195_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to195_input_global_id_0_0_stall_in_reg_195_NO_SHIFT_REG),
	.valid_out(rnode_4to195_input_global_id_0_0_valid_out_reg_195_NO_SHIFT_REG),
	.stall_out(rnode_4to195_input_global_id_0_0_stall_out_reg_195_NO_SHIFT_REG),
	.data_in(rnode_1to4_input_global_id_0_2_NO_SHIFT_REG),
	.data_out(rnode_4to195_input_global_id_0_0_reg_195_NO_SHIFT_REG)
);

defparam rnode_4to195_input_global_id_0_0_reg_195_fifo.DEPTH = 192;
defparam rnode_4to195_input_global_id_0_0_reg_195_fifo.DATA_WIDTH = 32;
defparam rnode_4to195_input_global_id_0_0_reg_195_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to195_input_global_id_0_0_reg_195_fifo.IMPL = "ram";

assign rnode_4to195_input_global_id_0_0_reg_195_inputs_ready_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_valid_out_2_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_stall_in_2_NO_SHIFT_REG = rnode_4to195_input_global_id_0_0_stall_out_reg_195_NO_SHIFT_REG;
assign rnode_4to195_input_global_id_0_0_NO_SHIFT_REG = rnode_4to195_input_global_id_0_0_reg_195_NO_SHIFT_REG;
assign rnode_4to195_input_global_id_0_0_stall_in_reg_195_NO_SHIFT_REG = rnode_4to195_input_global_id_0_0_stall_in_NO_SHIFT_REG;
assign rnode_4to195_input_global_id_0_0_valid_out_NO_SHIFT_REG = rnode_4to195_input_global_id_0_0_valid_out_reg_195_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_lftr_wideiv_valid_out_1;
wire local_bb2_lftr_wideiv_stall_in_1;
 reg local_bb2_lftr_wideiv_consumed_1_NO_SHIFT_REG;
wire local_bb2_exitcond_valid_out;
wire local_bb2_exitcond_stall_in;
 reg local_bb2_exitcond_consumed_0_NO_SHIFT_REG;
wire local_bb2_exitcond_inputs_ready;
wire local_bb2_exitcond_stall_local;
wire local_bb2_exitcond;

assign local_bb2_exitcond_inputs_ready = merge_node_valid_out_0_NO_SHIFT_REG;
assign local_bb2_exitcond = (local_bb2_lftr_wideiv == input_c1f2);
assign local_bb2_exitcond_stall_local = ((local_bb2_lftr_wideiv_stall_in_1 & ~(local_bb2_lftr_wideiv_consumed_1_NO_SHIFT_REG)) | (local_bb2_exitcond_stall_in & ~(local_bb2_exitcond_consumed_0_NO_SHIFT_REG)));
assign local_bb2_lftr_wideiv_valid_out_1 = (local_bb2_exitcond_inputs_ready & ~(local_bb2_lftr_wideiv_consumed_1_NO_SHIFT_REG));
assign local_bb2_exitcond_valid_out = (local_bb2_exitcond_inputs_ready & ~(local_bb2_exitcond_consumed_0_NO_SHIFT_REG));
assign merge_node_stall_in_0 = (|local_bb2_exitcond_stall_local);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_lftr_wideiv_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_exitcond_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_lftr_wideiv_consumed_1_NO_SHIFT_REG <= (local_bb2_exitcond_inputs_ready & (local_bb2_lftr_wideiv_consumed_1_NO_SHIFT_REG | ~(local_bb2_lftr_wideiv_stall_in_1)) & local_bb2_exitcond_stall_local);
		local_bb2_exitcond_consumed_0_NO_SHIFT_REG <= (local_bb2_exitcond_inputs_ready & (local_bb2_exitcond_consumed_0_NO_SHIFT_REG | ~(local_bb2_exitcond_stall_in)) & local_bb2_exitcond_stall_local);
	end
end


// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_4to4_bb2_mul4_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb2_mul4_0_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb2_mul4_0_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_4to4_bb2_mul4_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to4_bb2_mul4_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to4_bb2_mul4_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_4to4_bb2_mul4_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_4to4_bb2_mul4_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb2_mul4),
	.data_out(rnode_4to4_bb2_mul4_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_4to4_bb2_mul4_0_reg_4_fifo.DEPTH = 3;
defparam rnode_4to4_bb2_mul4_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_4to4_bb2_mul4_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to4_bb2_mul4_0_reg_4_fifo.IMPL = "zl_reg";

assign rnode_4to4_bb2_mul4_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb2_mul4_valid_out_NO_SHIFT_REG;
assign local_bb2_mul4_stall_in = rnode_4to4_bb2_mul4_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb2_mul4_0_NO_SHIFT_REG = rnode_4to4_bb2_mul4_0_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb2_mul4_0_stall_in_reg_4_NO_SHIFT_REG = rnode_4to4_bb2_mul4_0_stall_in_NO_SHIFT_REG;
assign rnode_4to4_bb2_mul4_0_valid_out_NO_SHIFT_REG = rnode_4to4_bb2_mul4_0_valid_out_reg_4_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_194to195_indvars_iv_0_valid_out_NO_SHIFT_REG;
 logic rnode_194to195_indvars_iv_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_194to195_indvars_iv_0_NO_SHIFT_REG;
 logic rnode_194to195_indvars_iv_0_reg_195_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_194to195_indvars_iv_0_reg_195_NO_SHIFT_REG;
 logic rnode_194to195_indvars_iv_0_valid_out_reg_195_NO_SHIFT_REG;
 logic rnode_194to195_indvars_iv_0_stall_in_reg_195_NO_SHIFT_REG;
 logic rnode_194to195_indvars_iv_0_stall_out_reg_195_NO_SHIFT_REG;

acl_data_fifo rnode_194to195_indvars_iv_0_reg_195_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_194to195_indvars_iv_0_reg_195_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_194to195_indvars_iv_0_stall_in_reg_195_NO_SHIFT_REG),
	.valid_out(rnode_194to195_indvars_iv_0_valid_out_reg_195_NO_SHIFT_REG),
	.stall_out(rnode_194to195_indvars_iv_0_stall_out_reg_195_NO_SHIFT_REG),
	.data_in(rnode_4to194_indvars_iv_0_NO_SHIFT_REG),
	.data_out(rnode_194to195_indvars_iv_0_reg_195_NO_SHIFT_REG)
);

defparam rnode_194to195_indvars_iv_0_reg_195_fifo.DEPTH = 2;
defparam rnode_194to195_indvars_iv_0_reg_195_fifo.DATA_WIDTH = 64;
defparam rnode_194to195_indvars_iv_0_reg_195_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_194to195_indvars_iv_0_reg_195_fifo.IMPL = "ll_reg";

assign rnode_194to195_indvars_iv_0_reg_195_inputs_ready_NO_SHIFT_REG = rnode_4to194_indvars_iv_0_valid_out_NO_SHIFT_REG;
assign rnode_4to194_indvars_iv_0_stall_in_NO_SHIFT_REG = rnode_194to195_indvars_iv_0_stall_out_reg_195_NO_SHIFT_REG;
assign rnode_194to195_indvars_iv_0_NO_SHIFT_REG = rnode_194to195_indvars_iv_0_reg_195_NO_SHIFT_REG;
assign rnode_194to195_indvars_iv_0_stall_in_reg_195_NO_SHIFT_REG = rnode_194to195_indvars_iv_0_stall_in_NO_SHIFT_REG;
assign rnode_194to195_indvars_iv_0_valid_out_NO_SHIFT_REG = rnode_194to195_indvars_iv_0_valid_out_reg_195_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb2_var__u0_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_4to5_bb2_var__u0_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_4to5_bb2_var__u0_0_NO_SHIFT_REG;
 logic rnode_4to5_bb2_var__u0_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_4to5_bb2_var__u0_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_4to5_bb2_var__u0_1_NO_SHIFT_REG;
 logic rnode_4to5_bb2_var__u0_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_4to5_bb2_var__u0_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_var__u0_0_valid_out_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_var__u0_0_stall_in_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_var__u0_0_stall_out_reg_5_NO_SHIFT_REG;
 logic [63:0] rnode_4to5_bb2_var__u0_0_reg_5_NO_SHIFT_REG_fa;

acl_multi_fanout_adaptor rnode_4to5_bb2_var__u0_0_reg_5_fanout_adaptor (
	.clock(clock),
	.resetn(resetn),
	.data_in(rnode_4to5_bb2_var__u0_0_reg_5_NO_SHIFT_REG),
	.valid_in(rnode_4to5_bb2_var__u0_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb2_var__u0_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.data_out(rnode_4to5_bb2_var__u0_0_reg_5_NO_SHIFT_REG_fa),
	.valid_out({rnode_4to5_bb2_var__u0_0_valid_out_0_NO_SHIFT_REG, rnode_4to5_bb2_var__u0_0_valid_out_1_NO_SHIFT_REG}),
	.stall_in({rnode_4to5_bb2_var__u0_0_stall_in_0_NO_SHIFT_REG, rnode_4to5_bb2_var__u0_0_stall_in_1_NO_SHIFT_REG})
);

defparam rnode_4to5_bb2_var__u0_0_reg_5_fanout_adaptor.DATA_WIDTH = 64;
defparam rnode_4to5_bb2_var__u0_0_reg_5_fanout_adaptor.NUM_FANOUTS = 2;

acl_data_fifo rnode_4to5_bb2_var__u0_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb2_var__u0_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb2_var__u0_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb2_var__u0_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb2_var__u0_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb2_var__u0),
	.data_out(rnode_4to5_bb2_var__u0_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb2_var__u0_0_reg_5_fifo.DEPTH = 2;
defparam rnode_4to5_bb2_var__u0_0_reg_5_fifo.DATA_WIDTH = 64;
defparam rnode_4to5_bb2_var__u0_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to5_bb2_var__u0_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_4to5_bb2_var__u0_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb2_var__u0_valid_out;
assign local_bb2_var__u0_stall_in = rnode_4to5_bb2_var__u0_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb2_var__u0_0_NO_SHIFT_REG = rnode_4to5_bb2_var__u0_0_reg_5_NO_SHIFT_REG_fa;
assign rnode_4to5_bb2_var__u0_1_NO_SHIFT_REG = rnode_4to5_bb2_var__u0_0_reg_5_NO_SHIFT_REG_fa;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_195to196_var__0_valid_out_NO_SHIFT_REG;
 logic rnode_195to196_var__0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_195to196_var__0_NO_SHIFT_REG;
 logic rnode_195to196_var__0_reg_196_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_195to196_var__0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_var__0_valid_out_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_var__0_stall_in_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_var__0_stall_out_reg_196_NO_SHIFT_REG;

acl_data_fifo rnode_195to196_var__0_reg_196_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_195to196_var__0_reg_196_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_195to196_var__0_stall_in_reg_196_NO_SHIFT_REG),
	.valid_out(rnode_195to196_var__0_valid_out_reg_196_NO_SHIFT_REG),
	.stall_out(rnode_195to196_var__0_stall_out_reg_196_NO_SHIFT_REG),
	.data_in(rnode_4to195_var__0_NO_SHIFT_REG),
	.data_out(rnode_195to196_var__0_reg_196_NO_SHIFT_REG)
);

defparam rnode_195to196_var__0_reg_196_fifo.DEPTH = 2;
defparam rnode_195to196_var__0_reg_196_fifo.DATA_WIDTH = 64;
defparam rnode_195to196_var__0_reg_196_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_195to196_var__0_reg_196_fifo.IMPL = "ll_reg";

assign rnode_195to196_var__0_reg_196_inputs_ready_NO_SHIFT_REG = rnode_4to195_var__0_valid_out_NO_SHIFT_REG;
assign rnode_4to195_var__0_stall_in_NO_SHIFT_REG = rnode_195to196_var__0_stall_out_reg_196_NO_SHIFT_REG;
assign rnode_195to196_var__0_NO_SHIFT_REG = rnode_195to196_var__0_reg_196_NO_SHIFT_REG;
assign rnode_195to196_var__0_stall_in_reg_196_NO_SHIFT_REG = rnode_195to196_var__0_stall_in_NO_SHIFT_REG;
assign rnode_195to196_var__0_valid_out_NO_SHIFT_REG = rnode_195to196_var__0_valid_out_reg_196_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_195to196_input_global_id_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_0_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_195to196_input_global_id_0_0_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_0_0_reg_196_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_195to196_input_global_id_0_0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_0_0_valid_out_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_0_0_stall_in_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_input_global_id_0_0_stall_out_reg_196_NO_SHIFT_REG;

acl_data_fifo rnode_195to196_input_global_id_0_0_reg_196_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_195to196_input_global_id_0_0_reg_196_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_195to196_input_global_id_0_0_stall_in_reg_196_NO_SHIFT_REG),
	.valid_out(rnode_195to196_input_global_id_0_0_valid_out_reg_196_NO_SHIFT_REG),
	.stall_out(rnode_195to196_input_global_id_0_0_stall_out_reg_196_NO_SHIFT_REG),
	.data_in(rnode_4to195_input_global_id_0_0_NO_SHIFT_REG),
	.data_out(rnode_195to196_input_global_id_0_0_reg_196_NO_SHIFT_REG)
);

defparam rnode_195to196_input_global_id_0_0_reg_196_fifo.DEPTH = 2;
defparam rnode_195to196_input_global_id_0_0_reg_196_fifo.DATA_WIDTH = 32;
defparam rnode_195to196_input_global_id_0_0_reg_196_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_195to196_input_global_id_0_0_reg_196_fifo.IMPL = "ll_reg";

assign rnode_195to196_input_global_id_0_0_reg_196_inputs_ready_NO_SHIFT_REG = rnode_4to195_input_global_id_0_0_valid_out_NO_SHIFT_REG;
assign rnode_4to195_input_global_id_0_0_stall_in_NO_SHIFT_REG = rnode_195to196_input_global_id_0_0_stall_out_reg_196_NO_SHIFT_REG;
assign rnode_195to196_input_global_id_0_0_NO_SHIFT_REG = rnode_195to196_input_global_id_0_0_reg_196_NO_SHIFT_REG;
assign rnode_195to196_input_global_id_0_0_stall_in_reg_196_NO_SHIFT_REG = rnode_195to196_input_global_id_0_0_stall_in_NO_SHIFT_REG;
assign rnode_195to196_input_global_id_0_0_valid_out_NO_SHIFT_REG = rnode_195to196_input_global_id_0_0_valid_out_reg_196_NO_SHIFT_REG;

// This section implements a registered operation.
// 
wire local_bb2_mul4_1_inputs_ready;
 reg local_bb2_mul4_1_valid_out_NO_SHIFT_REG;
wire local_bb2_mul4_1_stall_in;
wire local_bb2_mul4_1_output_regs_ready;
wire [31:0] local_bb2_mul4_1;
 reg local_bb2_mul4_1_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul4_1_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul4_1_causedstall;

acl_int_mult32s_s5 int_module_local_bb2_mul4_1 (
	.clock(clock),
	.dataa(local_bb2_lftr_wideiv),
	.datab(input_col_m2),
	.enable(local_bb2_mul4_1_output_regs_ready),
	.result(local_bb2_mul4_1)
);

defparam int_module_local_bb2_mul4_1.INPUT1_WIDTH = 32;
defparam int_module_local_bb2_mul4_1.INPUT2_WIDTH = 32;

assign local_bb2_mul4_1_inputs_ready = local_bb2_lftr_wideiv_valid_out_1;
assign local_bb2_mul4_1_output_regs_ready = (&(~(local_bb2_mul4_1_valid_out_NO_SHIFT_REG) | ~(local_bb2_mul4_1_stall_in)));
assign local_bb2_lftr_wideiv_stall_in_1 = (~(local_bb2_mul4_1_output_regs_ready) | ~(local_bb2_mul4_1_inputs_ready));
assign local_bb2_mul4_1_causedstall = (local_bb2_mul4_1_inputs_ready && (~(local_bb2_mul4_1_output_regs_ready) && !(~(local_bb2_mul4_1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul4_1_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul4_1_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul4_1_output_regs_ready)
		begin
			local_bb2_mul4_1_valid_pipe_0_NO_SHIFT_REG <= local_bb2_mul4_1_inputs_ready;
			local_bb2_mul4_1_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul4_1_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul4_1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul4_1_output_regs_ready)
		begin
			local_bb2_mul4_1_valid_out_NO_SHIFT_REG <= local_bb2_mul4_1_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb2_mul4_1_stall_in))
			begin
				local_bb2_mul4_1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_1to5_bb2_exitcond_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_1_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_valid_out_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_stall_in_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_stall_out_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb2_exitcond_0_reg_5_NO_SHIFT_REG_fa;

acl_multi_fanout_adaptor rnode_1to5_bb2_exitcond_0_reg_5_fanout_adaptor (
	.clock(clock),
	.resetn(resetn),
	.data_in(rnode_1to5_bb2_exitcond_0_reg_5_NO_SHIFT_REG),
	.valid_in(rnode_1to5_bb2_exitcond_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_1to5_bb2_exitcond_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.data_out(rnode_1to5_bb2_exitcond_0_reg_5_NO_SHIFT_REG_fa),
	.valid_out({rnode_1to5_bb2_exitcond_0_valid_out_0_NO_SHIFT_REG, rnode_1to5_bb2_exitcond_0_valid_out_1_NO_SHIFT_REG}),
	.stall_in({rnode_1to5_bb2_exitcond_0_stall_in_0_NO_SHIFT_REG, rnode_1to5_bb2_exitcond_0_stall_in_1_NO_SHIFT_REG})
);

defparam rnode_1to5_bb2_exitcond_0_reg_5_fanout_adaptor.DATA_WIDTH = 1;
defparam rnode_1to5_bb2_exitcond_0_reg_5_fanout_adaptor.NUM_FANOUTS = 2;

acl_data_fifo rnode_1to5_bb2_exitcond_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to5_bb2_exitcond_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to5_bb2_exitcond_0_stall_in_0_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_1to5_bb2_exitcond_0_valid_out_0_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_1to5_bb2_exitcond_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb2_exitcond),
	.data_out(rnode_1to5_bb2_exitcond_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_1to5_bb2_exitcond_0_reg_5_fifo.DEPTH = 5;
defparam rnode_1to5_bb2_exitcond_0_reg_5_fifo.DATA_WIDTH = 1;
defparam rnode_1to5_bb2_exitcond_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to5_bb2_exitcond_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_1to5_bb2_exitcond_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb2_exitcond_valid_out;
assign local_bb2_exitcond_stall_in = rnode_1to5_bb2_exitcond_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_1to5_bb2_exitcond_0_NO_SHIFT_REG = rnode_1to5_bb2_exitcond_0_reg_5_NO_SHIFT_REG_fa;
assign rnode_1to5_bb2_exitcond_1_NO_SHIFT_REG = rnode_1to5_bb2_exitcond_0_reg_5_NO_SHIFT_REG_fa;

// This section implements an unregistered operation.
// 
wire local_bb2_add5_valid_out;
wire local_bb2_add5_stall_in;
wire local_bb2_add5_inputs_ready;
wire local_bb2_add5_stall_local;
wire [31:0] local_bb2_add5;

assign local_bb2_add5_inputs_ready = (rnode_1to4_input_global_id_0_0_valid_out_0_NO_SHIFT_REG & rnode_4to4_bb2_mul4_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add5 = (rnode_4to4_bb2_mul4_0_NO_SHIFT_REG + rnode_1to4_input_global_id_0_0_NO_SHIFT_REG);
assign local_bb2_add5_valid_out = local_bb2_add5_inputs_ready;
assign local_bb2_add5_stall_local = local_bb2_add5_stall_in;
assign rnode_1to4_input_global_id_0_0_stall_in_0_NO_SHIFT_REG = (local_bb2_add5_stall_local | ~(local_bb2_add5_inputs_ready));
assign rnode_4to4_bb2_mul4_0_stall_in_NO_SHIFT_REG = (local_bb2_add5_stall_local | ~(local_bb2_add5_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb2_indvars_iv_next_1_valid_out;
wire local_bb2_indvars_iv_next_1_stall_in;
wire local_bb2_indvars_iv_next_1_inputs_ready;
wire local_bb2_indvars_iv_next_1_stall_local;
wire [63:0] local_bb2_indvars_iv_next_1;

assign local_bb2_indvars_iv_next_1_inputs_ready = rnode_194to195_indvars_iv_0_valid_out_NO_SHIFT_REG;
assign local_bb2_indvars_iv_next_1 = (rnode_194to195_indvars_iv_0_NO_SHIFT_REG + 64'h2);
assign local_bb2_indvars_iv_next_1_valid_out = local_bb2_indvars_iv_next_1_inputs_ready;
assign local_bb2_indvars_iv_next_1_stall_local = local_bb2_indvars_iv_next_1_stall_in;
assign rnode_194to195_indvars_iv_0_stall_in_NO_SHIFT_REG = (|local_bb2_indvars_iv_next_1_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx_stall_local;
wire [63:0] local_bb2_arrayidx;

assign local_bb2_arrayidx = (input_m1r + (rnode_4to5_bb2_var__u0_0_NO_SHIFT_REG << 6'h2));

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx12_stall_local;
wire [63:0] local_bb2_arrayidx12;

assign local_bb2_arrayidx12 = (input_m1i + (rnode_4to5_bb2_var__u0_1_NO_SHIFT_REG << 6'h2));

// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_4to4_bb2_mul4_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb2_mul4_1_0_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_1_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb2_mul4_1_0_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_1_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_1_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb2_mul4_1_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_4to4_bb2_mul4_1_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to4_bb2_mul4_1_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to4_bb2_mul4_1_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_4to4_bb2_mul4_1_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_4to4_bb2_mul4_1_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb2_mul4_1),
	.data_out(rnode_4to4_bb2_mul4_1_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_4to4_bb2_mul4_1_0_reg_4_fifo.DEPTH = 3;
defparam rnode_4to4_bb2_mul4_1_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_4to4_bb2_mul4_1_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to4_bb2_mul4_1_0_reg_4_fifo.IMPL = "zl_reg";

assign rnode_4to4_bb2_mul4_1_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb2_mul4_1_valid_out_NO_SHIFT_REG;
assign local_bb2_mul4_1_stall_in = rnode_4to4_bb2_mul4_1_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb2_mul4_1_0_NO_SHIFT_REG = rnode_4to4_bb2_mul4_1_0_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb2_mul4_1_0_stall_in_reg_4_NO_SHIFT_REG = rnode_4to4_bb2_mul4_1_0_stall_in_NO_SHIFT_REG;
assign rnode_4to4_bb2_mul4_1_0_valid_out_NO_SHIFT_REG = rnode_4to4_bb2_mul4_1_0_valid_out_reg_4_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp3_NEG_or49_valid_out;
wire local_bb2_cmp3_NEG_or49_stall_in;
wire local_bb2_cmp3_NEG_or49_inputs_ready;
wire local_bb2_cmp3_NEG_or49_stall_local;
wire local_bb2_cmp3_NEG_or49;

assign local_bb2_cmp3_NEG_or49_inputs_ready = rnode_1to5_bb2_exitcond_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_cmp3_NEG_or49 = (rnode_1to5_bb2_exitcond_0_NO_SHIFT_REG | input_wii_cmp3_NEG);
assign local_bb2_cmp3_NEG_or49_valid_out = local_bb2_cmp3_NEG_or49_inputs_ready;
assign local_bb2_cmp3_NEG_or49_stall_local = local_bb2_cmp3_NEG_or49_stall_in;
assign rnode_1to5_bb2_exitcond_0_stall_in_0_NO_SHIFT_REG = (|local_bb2_cmp3_NEG_or49_stall_local);

// Register node:
//  * latency = 190
//  * capacity = 190
 logic rnode_5to195_bb2_exitcond_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to195_bb2_exitcond_0_stall_in_NO_SHIFT_REG;
 logic rnode_5to195_bb2_exitcond_0_NO_SHIFT_REG;
 logic rnode_5to195_bb2_exitcond_0_reg_195_inputs_ready_NO_SHIFT_REG;
 logic rnode_5to195_bb2_exitcond_0_reg_195_NO_SHIFT_REG;
 logic rnode_5to195_bb2_exitcond_0_valid_out_reg_195_NO_SHIFT_REG;
 logic rnode_5to195_bb2_exitcond_0_stall_in_reg_195_NO_SHIFT_REG;
 logic rnode_5to195_bb2_exitcond_0_stall_out_reg_195_NO_SHIFT_REG;

acl_data_fifo rnode_5to195_bb2_exitcond_0_reg_195_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to195_bb2_exitcond_0_reg_195_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to195_bb2_exitcond_0_stall_in_reg_195_NO_SHIFT_REG),
	.valid_out(rnode_5to195_bb2_exitcond_0_valid_out_reg_195_NO_SHIFT_REG),
	.stall_out(rnode_5to195_bb2_exitcond_0_stall_out_reg_195_NO_SHIFT_REG),
	.data_in(rnode_1to5_bb2_exitcond_1_NO_SHIFT_REG),
	.data_out(rnode_5to195_bb2_exitcond_0_reg_195_NO_SHIFT_REG)
);

defparam rnode_5to195_bb2_exitcond_0_reg_195_fifo.DEPTH = 191;
defparam rnode_5to195_bb2_exitcond_0_reg_195_fifo.DATA_WIDTH = 1;
defparam rnode_5to195_bb2_exitcond_0_reg_195_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_5to195_bb2_exitcond_0_reg_195_fifo.IMPL = "ram";

assign rnode_5to195_bb2_exitcond_0_reg_195_inputs_ready_NO_SHIFT_REG = rnode_1to5_bb2_exitcond_0_valid_out_1_NO_SHIFT_REG;
assign rnode_1to5_bb2_exitcond_0_stall_in_1_NO_SHIFT_REG = rnode_5to195_bb2_exitcond_0_stall_out_reg_195_NO_SHIFT_REG;
assign rnode_5to195_bb2_exitcond_0_NO_SHIFT_REG = rnode_5to195_bb2_exitcond_0_reg_195_NO_SHIFT_REG;
assign rnode_5to195_bb2_exitcond_0_stall_in_reg_195_NO_SHIFT_REG = rnode_5to195_bb2_exitcond_0_stall_in_NO_SHIFT_REG;
assign rnode_5to195_bb2_exitcond_0_valid_out_NO_SHIFT_REG = rnode_5to195_bb2_exitcond_0_valid_out_reg_195_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb2_add5_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb2_add5_0_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb2_add5_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb2_add5_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb2_add5_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb2_add5_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb2_add5_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb2_add5_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb2_add5),
	.data_out(rnode_4to5_bb2_add5_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb2_add5_0_reg_5_fifo.DEPTH = 2;
defparam rnode_4to5_bb2_add5_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb2_add5_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to5_bb2_add5_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_4to5_bb2_add5_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb2_add5_valid_out;
assign local_bb2_add5_stall_in = rnode_4to5_bb2_add5_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb2_add5_0_NO_SHIFT_REG = rnode_4to5_bb2_add5_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb2_add5_0_stall_in_reg_5_NO_SHIFT_REG = rnode_4to5_bb2_add5_0_stall_in_NO_SHIFT_REG;
assign rnode_4to5_bb2_add5_0_valid_out_NO_SHIFT_REG = rnode_4to5_bb2_add5_0_valid_out_reg_5_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_0_NO_SHIFT_REG;
 logic [63:0] rnode_195to196_bb2_indvars_iv_next_1_0_NO_SHIFT_REG;
 logic rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_1_NO_SHIFT_REG;
 logic [63:0] rnode_195to196_bb2_indvars_iv_next_1_1_NO_SHIFT_REG;
 logic rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_bb2_indvars_iv_next_1_0_stall_out_reg_196_NO_SHIFT_REG;
 logic [63:0] rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_NO_SHIFT_REG_fa;

acl_multi_fanout_adaptor rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_fanout_adaptor (
	.clock(clock),
	.resetn(resetn),
	.data_in(rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_NO_SHIFT_REG),
	.valid_in(rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_0_reg_196_NO_SHIFT_REG),
	.stall_out(rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_0_reg_196_NO_SHIFT_REG),
	.data_out(rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_NO_SHIFT_REG_fa),
	.valid_out({rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_0_NO_SHIFT_REG, rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_1_NO_SHIFT_REG}),
	.stall_in({rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_0_NO_SHIFT_REG, rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_1_NO_SHIFT_REG})
);

defparam rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_fanout_adaptor.DATA_WIDTH = 64;
defparam rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_fanout_adaptor.NUM_FANOUTS = 2;

acl_data_fifo rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_0_reg_196_NO_SHIFT_REG),
	.valid_out(rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_0_reg_196_NO_SHIFT_REG),
	.stall_out(rnode_195to196_bb2_indvars_iv_next_1_0_stall_out_reg_196_NO_SHIFT_REG),
	.data_in(local_bb2_indvars_iv_next_1),
	.data_out(rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_NO_SHIFT_REG)
);

defparam rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_fifo.DEPTH = 2;
defparam rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_fifo.DATA_WIDTH = 64;
defparam rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_fifo.IMPL = "ll_reg";

assign rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_inputs_ready_NO_SHIFT_REG = local_bb2_indvars_iv_next_1_valid_out;
assign local_bb2_indvars_iv_next_1_stall_in = rnode_195to196_bb2_indvars_iv_next_1_0_stall_out_reg_196_NO_SHIFT_REG;
assign rnode_195to196_bb2_indvars_iv_next_1_0_NO_SHIFT_REG = rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_NO_SHIFT_REG_fa;
assign rnode_195to196_bb2_indvars_iv_next_1_1_NO_SHIFT_REG = rnode_195to196_bb2_indvars_iv_next_1_0_reg_196_NO_SHIFT_REG_fa;

// This section implements an unregistered operation.
// 
wire local_bb2_memcoalesce_m1r_bitcast_0_valid_out;
wire local_bb2_memcoalesce_m1r_bitcast_0_stall_in;
wire local_bb2_memcoalesce_m1r_bitcast_0_inputs_ready;
wire local_bb2_memcoalesce_m1r_bitcast_0_stall_local;
wire [63:0] local_bb2_memcoalesce_m1r_bitcast_0;

assign local_bb2_memcoalesce_m1r_bitcast_0_inputs_ready = rnode_4to5_bb2_var__u0_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_memcoalesce_m1r_bitcast_0 = local_bb2_arrayidx;
assign local_bb2_memcoalesce_m1r_bitcast_0_valid_out = local_bb2_memcoalesce_m1r_bitcast_0_inputs_ready;
assign local_bb2_memcoalesce_m1r_bitcast_0_stall_local = local_bb2_memcoalesce_m1r_bitcast_0_stall_in;
assign rnode_4to5_bb2_var__u0_0_stall_in_0_NO_SHIFT_REG = (|local_bb2_memcoalesce_m1r_bitcast_0_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb2_memcoalesce_m1i_bitcast_0_valid_out;
wire local_bb2_memcoalesce_m1i_bitcast_0_stall_in;
wire local_bb2_memcoalesce_m1i_bitcast_0_inputs_ready;
wire local_bb2_memcoalesce_m1i_bitcast_0_stall_local;
wire [63:0] local_bb2_memcoalesce_m1i_bitcast_0;

assign local_bb2_memcoalesce_m1i_bitcast_0_inputs_ready = rnode_4to5_bb2_var__u0_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_memcoalesce_m1i_bitcast_0 = local_bb2_arrayidx12;
assign local_bb2_memcoalesce_m1i_bitcast_0_valid_out = local_bb2_memcoalesce_m1i_bitcast_0_inputs_ready;
assign local_bb2_memcoalesce_m1i_bitcast_0_stall_local = local_bb2_memcoalesce_m1i_bitcast_0_stall_in;
assign rnode_4to5_bb2_var__u0_0_stall_in_1_NO_SHIFT_REG = (|local_bb2_memcoalesce_m1i_bitcast_0_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb2_add5_1_valid_out;
wire local_bb2_add5_1_stall_in;
wire local_bb2_add5_1_inputs_ready;
wire local_bb2_add5_1_stall_local;
wire [31:0] local_bb2_add5_1;

assign local_bb2_add5_1_inputs_ready = (rnode_1to4_input_global_id_0_0_valid_out_1_NO_SHIFT_REG & rnode_4to4_bb2_mul4_1_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add5_1 = (rnode_4to4_bb2_mul4_1_0_NO_SHIFT_REG + rnode_1to4_input_global_id_0_1_NO_SHIFT_REG);
assign local_bb2_add5_1_valid_out = local_bb2_add5_1_inputs_ready;
assign local_bb2_add5_1_stall_local = local_bb2_add5_1_stall_in;
assign rnode_1to4_input_global_id_0_0_stall_in_1_NO_SHIFT_REG = (local_bb2_add5_1_stall_local | ~(local_bb2_add5_1_inputs_ready));
assign rnode_4to4_bb2_mul4_1_0_stall_in_NO_SHIFT_REG = (local_bb2_add5_1_stall_local | ~(local_bb2_add5_1_inputs_ready));

// This section implements a staging register.
// 
wire rstag_5to5_bb2_cmp3_NEG_or49_valid_out_0;
wire rstag_5to5_bb2_cmp3_NEG_or49_stall_in_0;
 reg rstag_5to5_bb2_cmp3_NEG_or49_consumed_0_NO_SHIFT_REG;
wire rstag_5to5_bb2_cmp3_NEG_or49_valid_out_1;
wire rstag_5to5_bb2_cmp3_NEG_or49_stall_in_1;
 reg rstag_5to5_bb2_cmp3_NEG_or49_consumed_1_NO_SHIFT_REG;
wire rstag_5to5_bb2_cmp3_NEG_or49_inputs_ready;
wire rstag_5to5_bb2_cmp3_NEG_or49_stall_local;
 reg rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb2_cmp3_NEG_or49_combined_valid;
 reg rstag_5to5_bb2_cmp3_NEG_or49_staging_reg_NO_SHIFT_REG;
wire rstag_5to5_bb2_cmp3_NEG_or49;

assign rstag_5to5_bb2_cmp3_NEG_or49_inputs_ready = local_bb2_cmp3_NEG_or49_valid_out;
assign rstag_5to5_bb2_cmp3_NEG_or49 = (rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb2_cmp3_NEG_or49_staging_reg_NO_SHIFT_REG : local_bb2_cmp3_NEG_or49);
assign rstag_5to5_bb2_cmp3_NEG_or49_combined_valid = (rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG | rstag_5to5_bb2_cmp3_NEG_or49_inputs_ready);
assign rstag_5to5_bb2_cmp3_NEG_or49_stall_local = ((rstag_5to5_bb2_cmp3_NEG_or49_stall_in_0 & ~(rstag_5to5_bb2_cmp3_NEG_or49_consumed_0_NO_SHIFT_REG)) | (rstag_5to5_bb2_cmp3_NEG_or49_stall_in_1 & ~(rstag_5to5_bb2_cmp3_NEG_or49_consumed_1_NO_SHIFT_REG)));
assign rstag_5to5_bb2_cmp3_NEG_or49_valid_out_0 = (rstag_5to5_bb2_cmp3_NEG_or49_combined_valid & ~(rstag_5to5_bb2_cmp3_NEG_or49_consumed_0_NO_SHIFT_REG));
assign rstag_5to5_bb2_cmp3_NEG_or49_valid_out_1 = (rstag_5to5_bb2_cmp3_NEG_or49_combined_valid & ~(rstag_5to5_bb2_cmp3_NEG_or49_consumed_1_NO_SHIFT_REG));
assign local_bb2_cmp3_NEG_or49_stall_in = (|rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb2_cmp3_NEG_or49_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_5to5_bb2_cmp3_NEG_or49_stall_local)
		begin
			if (~(rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG))
			begin
				rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb2_cmp3_NEG_or49_inputs_ready;
			end
		end
		else
		begin
			rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_5to5_bb2_cmp3_NEG_or49_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb2_cmp3_NEG_or49_staging_reg_NO_SHIFT_REG <= local_bb2_cmp3_NEG_or49;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb2_cmp3_NEG_or49_consumed_0_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb2_cmp3_NEG_or49_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		rstag_5to5_bb2_cmp3_NEG_or49_consumed_0_NO_SHIFT_REG <= (rstag_5to5_bb2_cmp3_NEG_or49_combined_valid & (rstag_5to5_bb2_cmp3_NEG_or49_consumed_0_NO_SHIFT_REG | ~(rstag_5to5_bb2_cmp3_NEG_or49_stall_in_0)) & rstag_5to5_bb2_cmp3_NEG_or49_stall_local);
		rstag_5to5_bb2_cmp3_NEG_or49_consumed_1_NO_SHIFT_REG <= (rstag_5to5_bb2_cmp3_NEG_or49_combined_valid & (rstag_5to5_bb2_cmp3_NEG_or49_consumed_1_NO_SHIFT_REG | ~(rstag_5to5_bb2_cmp3_NEG_or49_stall_in_1)) & rstag_5to5_bb2_cmp3_NEG_or49_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_195to196_bb2_exitcond_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_1_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_reg_196_inputs_ready_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_valid_out_0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_stall_in_0_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_stall_out_reg_196_NO_SHIFT_REG;
 logic rnode_195to196_bb2_exitcond_0_reg_196_NO_SHIFT_REG_fa;

acl_multi_fanout_adaptor rnode_195to196_bb2_exitcond_0_reg_196_fanout_adaptor (
	.clock(clock),
	.resetn(resetn),
	.data_in(rnode_195to196_bb2_exitcond_0_reg_196_NO_SHIFT_REG),
	.valid_in(rnode_195to196_bb2_exitcond_0_valid_out_0_reg_196_NO_SHIFT_REG),
	.stall_out(rnode_195to196_bb2_exitcond_0_stall_in_0_reg_196_NO_SHIFT_REG),
	.data_out(rnode_195to196_bb2_exitcond_0_reg_196_NO_SHIFT_REG_fa),
	.valid_out({rnode_195to196_bb2_exitcond_0_valid_out_0_NO_SHIFT_REG, rnode_195to196_bb2_exitcond_0_valid_out_1_NO_SHIFT_REG}),
	.stall_in({rnode_195to196_bb2_exitcond_0_stall_in_0_NO_SHIFT_REG, rnode_195to196_bb2_exitcond_0_stall_in_1_NO_SHIFT_REG})
);

defparam rnode_195to196_bb2_exitcond_0_reg_196_fanout_adaptor.DATA_WIDTH = 1;
defparam rnode_195to196_bb2_exitcond_0_reg_196_fanout_adaptor.NUM_FANOUTS = 2;

acl_data_fifo rnode_195to196_bb2_exitcond_0_reg_196_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_195to196_bb2_exitcond_0_reg_196_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_195to196_bb2_exitcond_0_stall_in_0_reg_196_NO_SHIFT_REG),
	.valid_out(rnode_195to196_bb2_exitcond_0_valid_out_0_reg_196_NO_SHIFT_REG),
	.stall_out(rnode_195to196_bb2_exitcond_0_stall_out_reg_196_NO_SHIFT_REG),
	.data_in(rnode_5to195_bb2_exitcond_0_NO_SHIFT_REG),
	.data_out(rnode_195to196_bb2_exitcond_0_reg_196_NO_SHIFT_REG)
);

defparam rnode_195to196_bb2_exitcond_0_reg_196_fifo.DEPTH = 2;
defparam rnode_195to196_bb2_exitcond_0_reg_196_fifo.DATA_WIDTH = 1;
defparam rnode_195to196_bb2_exitcond_0_reg_196_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_195to196_bb2_exitcond_0_reg_196_fifo.IMPL = "ll_reg";

assign rnode_195to196_bb2_exitcond_0_reg_196_inputs_ready_NO_SHIFT_REG = rnode_5to195_bb2_exitcond_0_valid_out_NO_SHIFT_REG;
assign rnode_5to195_bb2_exitcond_0_stall_in_NO_SHIFT_REG = rnode_195to196_bb2_exitcond_0_stall_out_reg_196_NO_SHIFT_REG;
assign rnode_195to196_bb2_exitcond_0_NO_SHIFT_REG = rnode_195to196_bb2_exitcond_0_reg_196_NO_SHIFT_REG_fa;
assign rnode_195to196_bb2_exitcond_1_NO_SHIFT_REG = rnode_195to196_bb2_exitcond_0_reg_196_NO_SHIFT_REG_fa;

// This section implements an unregistered operation.
// 
wire local_bb2_idxprom6_stall_local;
wire [63:0] local_bb2_idxprom6;

assign local_bb2_idxprom6[32] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[33] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[34] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[35] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[36] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[37] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[38] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[39] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[40] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[41] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[42] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[43] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[44] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[45] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[46] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[47] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[48] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[49] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[50] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[51] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[52] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[53] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[54] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[55] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[56] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[57] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[58] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[59] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[60] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[61] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[62] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[63] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6[31:0] = rnode_4to5_bb2_add5_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_lftr_wideiv_1_stall_local;
wire [31:0] local_bb2_lftr_wideiv_1;

assign local_bb2_lftr_wideiv_1 = rnode_195to196_bb2_indvars_iv_next_1_0_NO_SHIFT_REG[31:0];

// This section implements a registered operation.
// 
wire local_bb2_ld_memcoalesce_m1r_load_0_inputs_ready;
 reg local_bb2_ld_memcoalesce_m1r_load_0_valid_out_NO_SHIFT_REG;
wire local_bb2_ld_memcoalesce_m1r_load_0_stall_in;
wire local_bb2_ld_memcoalesce_m1r_load_0_output_regs_ready;
wire local_bb2_ld_memcoalesce_m1r_load_0_fu_stall_out;
wire local_bb2_ld_memcoalesce_m1r_load_0_fu_valid_out;
wire [63:0] local_bb2_ld_memcoalesce_m1r_load_0_lsu_dataout;
 reg [63:0] local_bb2_ld_memcoalesce_m1r_load_0_NO_SHIFT_REG;
wire local_bb2_ld_memcoalesce_m1r_load_0_causedstall;

lsu_top lsu_local_bb2_ld_memcoalesce_m1r_load_0 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld_memcoalesce_m1r_load_0_fu_stall_out),
	.i_valid(local_bb2_ld_memcoalesce_m1r_load_0_inputs_ready),
	.i_address(local_bb2_memcoalesce_m1r_bitcast_0),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(input_wii_cmp3_NEG),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld_memcoalesce_m1r_load_0_output_regs_ready)),
	.o_valid(local_bb2_ld_memcoalesce_m1r_load_0_fu_valid_out),
	.o_readdata(local_bb2_ld_memcoalesce_m1r_load_0_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld_memcoalesce_m1r_load_0_active),
	.avm_address(avm_local_bb2_ld_memcoalesce_m1r_load_0_address),
	.avm_read(avm_local_bb2_ld_memcoalesce_m1r_load_0_read),
	.avm_readdata(avm_local_bb2_ld_memcoalesce_m1r_load_0_readdata),
	.avm_write(avm_local_bb2_ld_memcoalesce_m1r_load_0_write),
	.avm_writeack(avm_local_bb2_ld_memcoalesce_m1r_load_0_writeack),
	.avm_burstcount(avm_local_bb2_ld_memcoalesce_m1r_load_0_burstcount),
	.avm_writedata(avm_local_bb2_ld_memcoalesce_m1r_load_0_writedata),
	.avm_byteenable(avm_local_bb2_ld_memcoalesce_m1r_load_0_byteenable),
	.avm_waitrequest(avm_local_bb2_ld_memcoalesce_m1r_load_0_waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld_memcoalesce_m1r_load_0_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.AWIDTH = 30;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.WIDTH_BYTES = 8;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.MWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.WRITEDATAWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.READ = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.ATOMIC = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.WIDTH = 64;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.MWIDTH = 256;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.MEMORY_SIDE_MEM_LATENCY = 64;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.USECACHING = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.ADDRSPACE = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1r_load_0.STYLE = "BURST-NON-ALIGNED";

assign local_bb2_ld_memcoalesce_m1r_load_0_inputs_ready = (local_bb2_memcoalesce_m1r_bitcast_0_valid_out & rnode_1to5_cmp3_NEG_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_ld_memcoalesce_m1r_load_0_output_regs_ready = (&(~(local_bb2_ld_memcoalesce_m1r_load_0_valid_out_NO_SHIFT_REG) | ~(local_bb2_ld_memcoalesce_m1r_load_0_stall_in)));
assign local_bb2_memcoalesce_m1r_bitcast_0_stall_in = (local_bb2_ld_memcoalesce_m1r_load_0_fu_stall_out | ~(local_bb2_ld_memcoalesce_m1r_load_0_inputs_ready));
assign rnode_1to5_cmp3_NEG_0_stall_in_0_NO_SHIFT_REG = (local_bb2_ld_memcoalesce_m1r_load_0_fu_stall_out | ~(local_bb2_ld_memcoalesce_m1r_load_0_inputs_ready));
assign local_bb2_ld_memcoalesce_m1r_load_0_causedstall = (local_bb2_ld_memcoalesce_m1r_load_0_inputs_ready && (local_bb2_ld_memcoalesce_m1r_load_0_fu_stall_out && !(~(local_bb2_ld_memcoalesce_m1r_load_0_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld_memcoalesce_m1r_load_0_NO_SHIFT_REG <= 'x;
		local_bb2_ld_memcoalesce_m1r_load_0_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld_memcoalesce_m1r_load_0_output_regs_ready)
		begin
			local_bb2_ld_memcoalesce_m1r_load_0_NO_SHIFT_REG <= local_bb2_ld_memcoalesce_m1r_load_0_lsu_dataout;
			local_bb2_ld_memcoalesce_m1r_load_0_valid_out_NO_SHIFT_REG <= local_bb2_ld_memcoalesce_m1r_load_0_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld_memcoalesce_m1r_load_0_stall_in))
			begin
				local_bb2_ld_memcoalesce_m1r_load_0_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_ld_memcoalesce_m1i_load_0_inputs_ready;
 reg local_bb2_ld_memcoalesce_m1i_load_0_valid_out_NO_SHIFT_REG;
wire local_bb2_ld_memcoalesce_m1i_load_0_stall_in;
wire local_bb2_ld_memcoalesce_m1i_load_0_output_regs_ready;
wire local_bb2_ld_memcoalesce_m1i_load_0_fu_stall_out;
wire local_bb2_ld_memcoalesce_m1i_load_0_fu_valid_out;
wire [63:0] local_bb2_ld_memcoalesce_m1i_load_0_lsu_dataout;
 reg [63:0] local_bb2_ld_memcoalesce_m1i_load_0_NO_SHIFT_REG;
wire local_bb2_ld_memcoalesce_m1i_load_0_causedstall;

lsu_top lsu_local_bb2_ld_memcoalesce_m1i_load_0 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld_memcoalesce_m1i_load_0_fu_stall_out),
	.i_valid(local_bb2_ld_memcoalesce_m1i_load_0_inputs_ready),
	.i_address(local_bb2_memcoalesce_m1i_bitcast_0),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(input_wii_cmp3_NEG),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld_memcoalesce_m1i_load_0_output_regs_ready)),
	.o_valid(local_bb2_ld_memcoalesce_m1i_load_0_fu_valid_out),
	.o_readdata(local_bb2_ld_memcoalesce_m1i_load_0_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld_memcoalesce_m1i_load_0_active),
	.avm_address(avm_local_bb2_ld_memcoalesce_m1i_load_0_address),
	.avm_read(avm_local_bb2_ld_memcoalesce_m1i_load_0_read),
	.avm_readdata(avm_local_bb2_ld_memcoalesce_m1i_load_0_readdata),
	.avm_write(avm_local_bb2_ld_memcoalesce_m1i_load_0_write),
	.avm_writeack(avm_local_bb2_ld_memcoalesce_m1i_load_0_writeack),
	.avm_burstcount(avm_local_bb2_ld_memcoalesce_m1i_load_0_burstcount),
	.avm_writedata(avm_local_bb2_ld_memcoalesce_m1i_load_0_writedata),
	.avm_byteenable(avm_local_bb2_ld_memcoalesce_m1i_load_0_byteenable),
	.avm_waitrequest(avm_local_bb2_ld_memcoalesce_m1i_load_0_waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld_memcoalesce_m1i_load_0_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.AWIDTH = 30;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.WIDTH_BYTES = 8;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.MWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.WRITEDATAWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.READ = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.ATOMIC = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.WIDTH = 64;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.MWIDTH = 256;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.MEMORY_SIDE_MEM_LATENCY = 64;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.USECACHING = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.ADDRSPACE = 1;
defparam lsu_local_bb2_ld_memcoalesce_m1i_load_0.STYLE = "BURST-NON-ALIGNED";

assign local_bb2_ld_memcoalesce_m1i_load_0_inputs_ready = (local_bb2_memcoalesce_m1i_bitcast_0_valid_out & rnode_1to5_cmp3_NEG_0_valid_out_1_NO_SHIFT_REG);
assign local_bb2_ld_memcoalesce_m1i_load_0_output_regs_ready = (&(~(local_bb2_ld_memcoalesce_m1i_load_0_valid_out_NO_SHIFT_REG) | ~(local_bb2_ld_memcoalesce_m1i_load_0_stall_in)));
assign local_bb2_memcoalesce_m1i_bitcast_0_stall_in = (local_bb2_ld_memcoalesce_m1i_load_0_fu_stall_out | ~(local_bb2_ld_memcoalesce_m1i_load_0_inputs_ready));
assign rnode_1to5_cmp3_NEG_0_stall_in_1_NO_SHIFT_REG = (local_bb2_ld_memcoalesce_m1i_load_0_fu_stall_out | ~(local_bb2_ld_memcoalesce_m1i_load_0_inputs_ready));
assign local_bb2_ld_memcoalesce_m1i_load_0_causedstall = (local_bb2_ld_memcoalesce_m1i_load_0_inputs_ready && (local_bb2_ld_memcoalesce_m1i_load_0_fu_stall_out && !(~(local_bb2_ld_memcoalesce_m1i_load_0_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld_memcoalesce_m1i_load_0_NO_SHIFT_REG <= 'x;
		local_bb2_ld_memcoalesce_m1i_load_0_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld_memcoalesce_m1i_load_0_output_regs_ready)
		begin
			local_bb2_ld_memcoalesce_m1i_load_0_NO_SHIFT_REG <= local_bb2_ld_memcoalesce_m1i_load_0_lsu_dataout;
			local_bb2_ld_memcoalesce_m1i_load_0_valid_out_NO_SHIFT_REG <= local_bb2_ld_memcoalesce_m1i_load_0_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld_memcoalesce_m1i_load_0_stall_in))
			begin
				local_bb2_ld_memcoalesce_m1i_load_0_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb2_add5_1_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_1_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_1_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb2_add5_1_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_1_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_1_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb2_add5_1_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb2_add5_1_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb2_add5_1_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb2_add5_1_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb2_add5_1_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb2_add5_1_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb2_add5_1),
	.data_out(rnode_4to5_bb2_add5_1_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb2_add5_1_0_reg_5_fifo.DEPTH = 2;
defparam rnode_4to5_bb2_add5_1_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb2_add5_1_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to5_bb2_add5_1_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_4to5_bb2_add5_1_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb2_add5_1_valid_out;
assign local_bb2_add5_1_stall_in = rnode_4to5_bb2_add5_1_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG = rnode_4to5_bb2_add5_1_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb2_add5_1_0_stall_in_reg_5_NO_SHIFT_REG = rnode_4to5_bb2_add5_1_0_stall_in_NO_SHIFT_REG;
assign rnode_4to5_bb2_add5_1_0_valid_out_NO_SHIFT_REG = rnode_4to5_bb2_add5_1_0_valid_out_reg_5_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx7_stall_local;
wire [63:0] local_bb2_arrayidx7;

assign local_bb2_arrayidx7 = (input_m2r + (local_bb2_idxprom6 << 6'h2));

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx7_valid_out;
wire local_bb2_arrayidx7_stall_in;
 reg local_bb2_arrayidx7_consumed_0_NO_SHIFT_REG;
wire local_bb2_arrayidx16_valid_out;
wire local_bb2_arrayidx16_stall_in;
 reg local_bb2_arrayidx16_consumed_0_NO_SHIFT_REG;
wire local_bb2_arrayidx16_inputs_ready;
wire local_bb2_arrayidx16_stall_local;
wire [63:0] local_bb2_arrayidx16;

assign local_bb2_arrayidx16_inputs_ready = rnode_4to5_bb2_add5_0_valid_out_NO_SHIFT_REG;
assign local_bb2_arrayidx16 = (input_m2i + (local_bb2_idxprom6 << 6'h2));
assign local_bb2_arrayidx16_stall_local = ((local_bb2_arrayidx7_stall_in & ~(local_bb2_arrayidx7_consumed_0_NO_SHIFT_REG)) | (local_bb2_arrayidx16_stall_in & ~(local_bb2_arrayidx16_consumed_0_NO_SHIFT_REG)));
assign local_bb2_arrayidx7_valid_out = (local_bb2_arrayidx16_inputs_ready & ~(local_bb2_arrayidx7_consumed_0_NO_SHIFT_REG));
assign local_bb2_arrayidx16_valid_out = (local_bb2_arrayidx16_inputs_ready & ~(local_bb2_arrayidx16_consumed_0_NO_SHIFT_REG));
assign rnode_4to5_bb2_add5_0_stall_in_NO_SHIFT_REG = (|local_bb2_arrayidx16_stall_local);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_arrayidx7_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_arrayidx16_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_arrayidx7_consumed_0_NO_SHIFT_REG <= (local_bb2_arrayidx16_inputs_ready & (local_bb2_arrayidx7_consumed_0_NO_SHIFT_REG | ~(local_bb2_arrayidx7_stall_in)) & local_bb2_arrayidx16_stall_local);
		local_bb2_arrayidx16_consumed_0_NO_SHIFT_REG <= (local_bb2_arrayidx16_inputs_ready & (local_bb2_arrayidx16_consumed_0_NO_SHIFT_REG | ~(local_bb2_arrayidx16_stall_in)) & local_bb2_arrayidx16_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_exitcond_1_stall_local;
wire local_bb2_exitcond_1;

assign local_bb2_exitcond_1 = (local_bb2_lftr_wideiv_1 == input_c1f2);

// Register node:
//  * latency = 0
//  * capacity = 80
 logic rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(local_bb2_ld_memcoalesce_m1r_load_0_NO_SHIFT_REG),
	.data_out(rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_NO_SHIFT_REG)
);

defparam rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_fifo.DEPTH = 81;
defparam rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_fifo.DATA_WIDTH = 64;
defparam rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_fifo.IMPL = "zl_ram";

assign rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_inputs_ready_NO_SHIFT_REG = local_bb2_ld_memcoalesce_m1r_load_0_valid_out_NO_SHIFT_REG;
assign local_bb2_ld_memcoalesce_m1r_load_0_stall_in = rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_NO_SHIFT_REG = rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_reg_165_NO_SHIFT_REG;
assign rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_in_reg_165_NO_SHIFT_REG = rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_in_NO_SHIFT_REG;
assign rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_valid_out_NO_SHIFT_REG = rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_valid_out_reg_165_NO_SHIFT_REG;

// Register node:
//  * latency = 0
//  * capacity = 80
 logic rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_valid_out_reg_165_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_in_reg_165_NO_SHIFT_REG;
 logic rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_out_reg_165_NO_SHIFT_REG;

acl_data_fifo rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_in_reg_165_NO_SHIFT_REG),
	.valid_out(rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_valid_out_reg_165_NO_SHIFT_REG),
	.stall_out(rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_out_reg_165_NO_SHIFT_REG),
	.data_in(local_bb2_ld_memcoalesce_m1i_load_0_NO_SHIFT_REG),
	.data_out(rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_NO_SHIFT_REG)
);

defparam rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_fifo.DEPTH = 81;
defparam rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_fifo.DATA_WIDTH = 64;
defparam rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_fifo.IMPL = "zl_ram";

assign rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_inputs_ready_NO_SHIFT_REG = local_bb2_ld_memcoalesce_m1i_load_0_valid_out_NO_SHIFT_REG;
assign local_bb2_ld_memcoalesce_m1i_load_0_stall_in = rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_out_reg_165_NO_SHIFT_REG;
assign rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_NO_SHIFT_REG = rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_reg_165_NO_SHIFT_REG;
assign rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_in_reg_165_NO_SHIFT_REG = rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_in_NO_SHIFT_REG;
assign rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_valid_out_NO_SHIFT_REG = rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_valid_out_reg_165_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_idxprom6_1_stall_local;
wire [63:0] local_bb2_idxprom6_1;

assign local_bb2_idxprom6_1[32] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[33] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[34] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[35] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[36] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[37] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[38] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[39] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[40] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[41] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[42] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[43] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[44] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[45] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[46] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[47] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[48] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[49] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[50] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[51] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[52] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[53] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[54] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[55] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[56] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[57] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[58] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[59] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[60] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[61] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[62] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[63] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG[31];
assign local_bb2_idxprom6_1[31:0] = rnode_4to5_bb2_add5_1_0_NO_SHIFT_REG;

// This section implements a staging register.
// 
wire rstag_5to5_bb2_arrayidx7_valid_out;
wire rstag_5to5_bb2_arrayidx7_stall_in;
wire rstag_5to5_bb2_arrayidx7_inputs_ready;
wire rstag_5to5_bb2_arrayidx7_stall_local;
 reg rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb2_arrayidx7_combined_valid;
 reg [63:0] rstag_5to5_bb2_arrayidx7_staging_reg_NO_SHIFT_REG;
wire [63:0] rstag_5to5_bb2_arrayidx7;

assign rstag_5to5_bb2_arrayidx7_inputs_ready = local_bb2_arrayidx7_valid_out;
assign rstag_5to5_bb2_arrayidx7 = (rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb2_arrayidx7_staging_reg_NO_SHIFT_REG : local_bb2_arrayidx7);
assign rstag_5to5_bb2_arrayidx7_combined_valid = (rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG | rstag_5to5_bb2_arrayidx7_inputs_ready);
assign rstag_5to5_bb2_arrayidx7_valid_out = rstag_5to5_bb2_arrayidx7_combined_valid;
assign rstag_5to5_bb2_arrayidx7_stall_local = rstag_5to5_bb2_arrayidx7_stall_in;
assign local_bb2_arrayidx7_stall_in = (|rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb2_arrayidx7_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_5to5_bb2_arrayidx7_stall_local)
		begin
			if (~(rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG))
			begin
				rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb2_arrayidx7_inputs_ready;
			end
		end
		else
		begin
			rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_5to5_bb2_arrayidx7_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb2_arrayidx7_staging_reg_NO_SHIFT_REG <= local_bb2_arrayidx7;
		end
	end
end


// This section implements a staging register.
// 
wire rstag_5to5_bb2_arrayidx16_valid_out;
wire rstag_5to5_bb2_arrayidx16_stall_in;
wire rstag_5to5_bb2_arrayidx16_inputs_ready;
wire rstag_5to5_bb2_arrayidx16_stall_local;
 reg rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb2_arrayidx16_combined_valid;
 reg [63:0] rstag_5to5_bb2_arrayidx16_staging_reg_NO_SHIFT_REG;
wire [63:0] rstag_5to5_bb2_arrayidx16;

assign rstag_5to5_bb2_arrayidx16_inputs_ready = local_bb2_arrayidx16_valid_out;
assign rstag_5to5_bb2_arrayidx16 = (rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb2_arrayidx16_staging_reg_NO_SHIFT_REG : local_bb2_arrayidx16);
assign rstag_5to5_bb2_arrayidx16_combined_valid = (rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG | rstag_5to5_bb2_arrayidx16_inputs_ready);
assign rstag_5to5_bb2_arrayidx16_valid_out = rstag_5to5_bb2_arrayidx16_combined_valid;
assign rstag_5to5_bb2_arrayidx16_stall_local = rstag_5to5_bb2_arrayidx16_stall_in;
assign local_bb2_arrayidx16_stall_in = (|rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb2_arrayidx16_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_5to5_bb2_arrayidx16_stall_local)
		begin
			if (~(rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG))
			begin
				rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb2_arrayidx16_inputs_ready;
			end
		end
		else
		begin
			rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_5to5_bb2_arrayidx16_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb2_arrayidx16_staging_reg_NO_SHIFT_REG <= local_bb2_arrayidx16;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2__24_demorgan_stall_local;
wire local_bb2__24_demorgan;

assign local_bb2__24_demorgan = (rnode_195to196_bb2_exitcond_0_NO_SHIFT_REG | local_bb2_exitcond_1);

// This section implements an unregistered operation.
// 
wire local_bb2_c0_eni1_stall_local;
wire [351:0] local_bb2_c0_eni1;

assign local_bb2_c0_eni1[31:0] = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
assign local_bb2_c0_eni1[95:32] = rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_NO_SHIFT_REG;
assign local_bb2_c0_eni1[351:96] = 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx7_1_stall_local;
wire [63:0] local_bb2_arrayidx7_1;

assign local_bb2_arrayidx7_1 = (input_m2r + (local_bb2_idxprom6_1 << 6'h2));

// This section implements an unregistered operation.
// 
wire local_bb2_arrayidx7_1_valid_out;
wire local_bb2_arrayidx7_1_stall_in;
 reg local_bb2_arrayidx7_1_consumed_0_NO_SHIFT_REG;
wire local_bb2_arrayidx16_1_valid_out;
wire local_bb2_arrayidx16_1_stall_in;
 reg local_bb2_arrayidx16_1_consumed_0_NO_SHIFT_REG;
wire local_bb2_arrayidx16_1_inputs_ready;
wire local_bb2_arrayidx16_1_stall_local;
wire [63:0] local_bb2_arrayidx16_1;

assign local_bb2_arrayidx16_1_inputs_ready = rnode_4to5_bb2_add5_1_0_valid_out_NO_SHIFT_REG;
assign local_bb2_arrayidx16_1 = (input_m2i + (local_bb2_idxprom6_1 << 6'h2));
assign local_bb2_arrayidx16_1_stall_local = ((local_bb2_arrayidx7_1_stall_in & ~(local_bb2_arrayidx7_1_consumed_0_NO_SHIFT_REG)) | (local_bb2_arrayidx16_1_stall_in & ~(local_bb2_arrayidx16_1_consumed_0_NO_SHIFT_REG)));
assign local_bb2_arrayidx7_1_valid_out = (local_bb2_arrayidx16_1_inputs_ready & ~(local_bb2_arrayidx7_1_consumed_0_NO_SHIFT_REG));
assign local_bb2_arrayidx16_1_valid_out = (local_bb2_arrayidx16_1_inputs_ready & ~(local_bb2_arrayidx16_1_consumed_0_NO_SHIFT_REG));
assign rnode_4to5_bb2_add5_1_0_stall_in_NO_SHIFT_REG = (|local_bb2_arrayidx16_1_stall_local);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_arrayidx7_1_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_arrayidx16_1_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_arrayidx7_1_consumed_0_NO_SHIFT_REG <= (local_bb2_arrayidx16_1_inputs_ready & (local_bb2_arrayidx7_1_consumed_0_NO_SHIFT_REG | ~(local_bb2_arrayidx7_1_stall_in)) & local_bb2_arrayidx16_1_stall_local);
		local_bb2_arrayidx16_1_consumed_0_NO_SHIFT_REG <= (local_bb2_arrayidx16_1_inputs_ready & (local_bb2_arrayidx16_1_consumed_0_NO_SHIFT_REG | ~(local_bb2_arrayidx16_1_stall_in)) & local_bb2_arrayidx16_1_stall_local);
	end
end


// This section implements a registered operation.
// 
wire local_bb2_ld__inputs_ready;
 reg local_bb2_ld__valid_out_NO_SHIFT_REG;
wire local_bb2_ld__stall_in;
wire local_bb2_ld__output_regs_ready;
wire local_bb2_ld__fu_stall_out;
wire local_bb2_ld__fu_valid_out;
wire [31:0] local_bb2_ld__lsu_dataout;
 reg [31:0] local_bb2_ld__NO_SHIFT_REG;
wire local_bb2_ld__causedstall;

lsu_top lsu_local_bb2_ld_ (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld__fu_stall_out),
	.i_valid(local_bb2_ld__inputs_ready),
	.i_address(rstag_5to5_bb2_arrayidx7),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(input_wii_cmp3_NEG),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld__output_regs_ready)),
	.o_valid(local_bb2_ld__fu_valid_out),
	.o_readdata(local_bb2_ld__lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld__active),
	.avm_address(avm_local_bb2_ld__address),
	.avm_read(avm_local_bb2_ld__read),
	.avm_readdata(avm_local_bb2_ld__readdata),
	.avm_write(avm_local_bb2_ld__write),
	.avm_writeack(avm_local_bb2_ld__writeack),
	.avm_burstcount(avm_local_bb2_ld__burstcount),
	.avm_writedata(avm_local_bb2_ld__writedata),
	.avm_byteenable(avm_local_bb2_ld__byteenable),
	.avm_waitrequest(avm_local_bb2_ld__waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld__readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld_.AWIDTH = 30;
defparam lsu_local_bb2_ld_.WIDTH_BYTES = 4;
defparam lsu_local_bb2_ld_.MWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld_.WRITEDATAWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld_.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb2_ld_.READ = 1;
defparam lsu_local_bb2_ld_.ATOMIC = 0;
defparam lsu_local_bb2_ld_.WIDTH = 32;
defparam lsu_local_bb2_ld_.MWIDTH = 256;
defparam lsu_local_bb2_ld_.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld_.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld_.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld_.MEMORY_SIDE_MEM_LATENCY = 61;
defparam lsu_local_bb2_ld_.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld_.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld_.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld_.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld_.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld_.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld_.USECACHING = 1;
defparam lsu_local_bb2_ld_.CACHESIZE = 256;
defparam lsu_local_bb2_ld_.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld_.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld_.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld_.ADDRSPACE = 1;
defparam lsu_local_bb2_ld_.STYLE = "BURST-COALESCED";

assign local_bb2_ld__inputs_ready = (rnode_1to5_cmp3_NEG_0_valid_out_2_NO_SHIFT_REG & rstag_5to5_bb2_arrayidx7_valid_out);
assign local_bb2_ld__output_regs_ready = (&(~(local_bb2_ld__valid_out_NO_SHIFT_REG) | ~(local_bb2_ld__stall_in)));
assign rnode_1to5_cmp3_NEG_0_stall_in_2_NO_SHIFT_REG = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign rstag_5to5_bb2_arrayidx7_stall_in = (local_bb2_ld__fu_stall_out | ~(local_bb2_ld__inputs_ready));
assign local_bb2_ld__causedstall = (local_bb2_ld__inputs_ready && (local_bb2_ld__fu_stall_out && !(~(local_bb2_ld__output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld__NO_SHIFT_REG <= 'x;
		local_bb2_ld__valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld__output_regs_ready)
		begin
			local_bb2_ld__NO_SHIFT_REG <= local_bb2_ld__lsu_dataout;
			local_bb2_ld__valid_out_NO_SHIFT_REG <= local_bb2_ld__fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld__stall_in))
			begin
				local_bb2_ld__valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_ld__u1_inputs_ready;
 reg local_bb2_ld__u1_valid_out_NO_SHIFT_REG;
wire local_bb2_ld__u1_stall_in;
wire local_bb2_ld__u1_output_regs_ready;
wire local_bb2_ld__u1_fu_stall_out;
wire local_bb2_ld__u1_fu_valid_out;
wire [31:0] local_bb2_ld__u1_lsu_dataout;
 reg [31:0] local_bb2_ld__u1_NO_SHIFT_REG;
wire local_bb2_ld__u1_causedstall;

lsu_top lsu_local_bb2_ld__u1 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld__u1_fu_stall_out),
	.i_valid(local_bb2_ld__u1_inputs_ready),
	.i_address(rstag_5to5_bb2_arrayidx16),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(input_wii_cmp3_NEG),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld__u1_output_regs_ready)),
	.o_valid(local_bb2_ld__u1_fu_valid_out),
	.o_readdata(local_bb2_ld__u1_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld__u1_active),
	.avm_address(avm_local_bb2_ld__u1_address),
	.avm_read(avm_local_bb2_ld__u1_read),
	.avm_readdata(avm_local_bb2_ld__u1_readdata),
	.avm_write(avm_local_bb2_ld__u1_write),
	.avm_writeack(avm_local_bb2_ld__u1_writeack),
	.avm_burstcount(avm_local_bb2_ld__u1_burstcount),
	.avm_writedata(avm_local_bb2_ld__u1_writedata),
	.avm_byteenable(avm_local_bb2_ld__u1_byteenable),
	.avm_waitrequest(avm_local_bb2_ld__u1_waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld__u1_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld__u1.AWIDTH = 30;
defparam lsu_local_bb2_ld__u1.WIDTH_BYTES = 4;
defparam lsu_local_bb2_ld__u1.MWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld__u1.WRITEDATAWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld__u1.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb2_ld__u1.READ = 1;
defparam lsu_local_bb2_ld__u1.ATOMIC = 0;
defparam lsu_local_bb2_ld__u1.WIDTH = 32;
defparam lsu_local_bb2_ld__u1.MWIDTH = 256;
defparam lsu_local_bb2_ld__u1.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld__u1.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld__u1.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld__u1.MEMORY_SIDE_MEM_LATENCY = 61;
defparam lsu_local_bb2_ld__u1.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld__u1.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld__u1.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld__u1.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld__u1.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld__u1.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld__u1.USECACHING = 1;
defparam lsu_local_bb2_ld__u1.CACHESIZE = 256;
defparam lsu_local_bb2_ld__u1.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld__u1.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld__u1.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld__u1.ADDRSPACE = 1;
defparam lsu_local_bb2_ld__u1.STYLE = "BURST-COALESCED";

assign local_bb2_ld__u1_inputs_ready = (rnode_1to5_cmp3_NEG_0_valid_out_3_NO_SHIFT_REG & rstag_5to5_bb2_arrayidx16_valid_out);
assign local_bb2_ld__u1_output_regs_ready = (&(~(local_bb2_ld__u1_valid_out_NO_SHIFT_REG) | ~(local_bb2_ld__u1_stall_in)));
assign rnode_1to5_cmp3_NEG_0_stall_in_3_NO_SHIFT_REG = (local_bb2_ld__u1_fu_stall_out | ~(local_bb2_ld__u1_inputs_ready));
assign rstag_5to5_bb2_arrayidx16_stall_in = (local_bb2_ld__u1_fu_stall_out | ~(local_bb2_ld__u1_inputs_ready));
assign local_bb2_ld__u1_causedstall = (local_bb2_ld__u1_inputs_ready && (local_bb2_ld__u1_fu_stall_out && !(~(local_bb2_ld__u1_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld__u1_NO_SHIFT_REG <= 'x;
		local_bb2_ld__u1_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld__u1_output_regs_ready)
		begin
			local_bb2_ld__u1_NO_SHIFT_REG <= local_bb2_ld__u1_lsu_dataout;
			local_bb2_ld__u1_valid_out_NO_SHIFT_REG <= local_bb2_ld__u1_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld__u1_stall_in))
			begin
				local_bb2_ld__u1_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2__24_demorgan_GUARD_valid_out;
wire local_bb2__24_demorgan_GUARD_stall_in;
wire local_bb2__24_demorgan_GUARD_inputs_ready;
wire local_bb2__24_demorgan_GUARD_stall_local;
wire local_bb2__24_demorgan_GUARD;

assign local_bb2__24_demorgan_GUARD_inputs_ready = (rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_0_NO_SHIFT_REG & rnode_195to196_bb2_exitcond_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2__24_demorgan_GUARD = (local_bb2__24_demorgan | input_wii_cmp3_NEG);
assign local_bb2__24_demorgan_GUARD_valid_out = local_bb2__24_demorgan_GUARD_inputs_ready;
assign local_bb2__24_demorgan_GUARD_stall_local = local_bb2__24_demorgan_GUARD_stall_in;
assign rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_0_NO_SHIFT_REG = (local_bb2__24_demorgan_GUARD_stall_local | ~(local_bb2__24_demorgan_GUARD_inputs_ready));
assign rnode_195to196_bb2_exitcond_0_stall_in_0_NO_SHIFT_REG = (local_bb2__24_demorgan_GUARD_stall_local | ~(local_bb2__24_demorgan_GUARD_inputs_ready));

// This section implements a staging register.
// 
wire rstag_5to5_bb2_arrayidx7_1_valid_out;
wire rstag_5to5_bb2_arrayidx7_1_stall_in;
wire rstag_5to5_bb2_arrayidx7_1_inputs_ready;
wire rstag_5to5_bb2_arrayidx7_1_stall_local;
 reg rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb2_arrayidx7_1_combined_valid;
 reg [63:0] rstag_5to5_bb2_arrayidx7_1_staging_reg_NO_SHIFT_REG;
wire [63:0] rstag_5to5_bb2_arrayidx7_1;

assign rstag_5to5_bb2_arrayidx7_1_inputs_ready = local_bb2_arrayidx7_1_valid_out;
assign rstag_5to5_bb2_arrayidx7_1 = (rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb2_arrayidx7_1_staging_reg_NO_SHIFT_REG : local_bb2_arrayidx7_1);
assign rstag_5to5_bb2_arrayidx7_1_combined_valid = (rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG | rstag_5to5_bb2_arrayidx7_1_inputs_ready);
assign rstag_5to5_bb2_arrayidx7_1_valid_out = rstag_5to5_bb2_arrayidx7_1_combined_valid;
assign rstag_5to5_bb2_arrayidx7_1_stall_local = rstag_5to5_bb2_arrayidx7_1_stall_in;
assign local_bb2_arrayidx7_1_stall_in = (|rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb2_arrayidx7_1_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_5to5_bb2_arrayidx7_1_stall_local)
		begin
			if (~(rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG))
			begin
				rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb2_arrayidx7_1_inputs_ready;
			end
		end
		else
		begin
			rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_5to5_bb2_arrayidx7_1_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb2_arrayidx7_1_staging_reg_NO_SHIFT_REG <= local_bb2_arrayidx7_1;
		end
	end
end


// This section implements a staging register.
// 
wire rstag_5to5_bb2_arrayidx16_1_valid_out;
wire rstag_5to5_bb2_arrayidx16_1_stall_in;
wire rstag_5to5_bb2_arrayidx16_1_inputs_ready;
wire rstag_5to5_bb2_arrayidx16_1_stall_local;
 reg rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb2_arrayidx16_1_combined_valid;
 reg [63:0] rstag_5to5_bb2_arrayidx16_1_staging_reg_NO_SHIFT_REG;
wire [63:0] rstag_5to5_bb2_arrayidx16_1;

assign rstag_5to5_bb2_arrayidx16_1_inputs_ready = local_bb2_arrayidx16_1_valid_out;
assign rstag_5to5_bb2_arrayidx16_1 = (rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb2_arrayidx16_1_staging_reg_NO_SHIFT_REG : local_bb2_arrayidx16_1);
assign rstag_5to5_bb2_arrayidx16_1_combined_valid = (rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG | rstag_5to5_bb2_arrayidx16_1_inputs_ready);
assign rstag_5to5_bb2_arrayidx16_1_valid_out = rstag_5to5_bb2_arrayidx16_1_combined_valid;
assign rstag_5to5_bb2_arrayidx16_1_stall_local = rstag_5to5_bb2_arrayidx16_1_stall_in;
assign local_bb2_arrayidx16_1_stall_in = (|rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb2_arrayidx16_1_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_5to5_bb2_arrayidx16_1_stall_local)
		begin
			if (~(rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG))
			begin
				rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb2_arrayidx16_1_inputs_ready;
			end
		end
		else
		begin
			rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_5to5_bb2_arrayidx16_1_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb2_arrayidx16_1_staging_reg_NO_SHIFT_REG <= local_bb2_arrayidx16_1;
		end
	end
end


// This section implements a staging register.
// 
wire rstag_165to165_bb2_ld__valid_out;
wire rstag_165to165_bb2_ld__stall_in;
wire rstag_165to165_bb2_ld__inputs_ready;
wire rstag_165to165_bb2_ld__stall_local;
 reg rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG;
wire rstag_165to165_bb2_ld__combined_valid;
 reg [31:0] rstag_165to165_bb2_ld__staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_165to165_bb2_ld_;

assign rstag_165to165_bb2_ld__inputs_ready = local_bb2_ld__valid_out_NO_SHIFT_REG;
assign rstag_165to165_bb2_ld_ = (rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG ? rstag_165to165_bb2_ld__staging_reg_NO_SHIFT_REG : local_bb2_ld__NO_SHIFT_REG);
assign rstag_165to165_bb2_ld__combined_valid = (rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG | rstag_165to165_bb2_ld__inputs_ready);
assign rstag_165to165_bb2_ld__valid_out = rstag_165to165_bb2_ld__combined_valid;
assign rstag_165to165_bb2_ld__stall_local = rstag_165to165_bb2_ld__stall_in;
assign local_bb2_ld__stall_in = (|rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_165to165_bb2_ld__staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_165to165_bb2_ld__stall_local)
		begin
			if (~(rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG))
			begin
				rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG <= rstag_165to165_bb2_ld__inputs_ready;
			end
		end
		else
		begin
			rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_165to165_bb2_ld__staging_valid_NO_SHIFT_REG))
		begin
			rstag_165to165_bb2_ld__staging_reg_NO_SHIFT_REG <= local_bb2_ld__NO_SHIFT_REG;
		end
	end
end


// This section implements a staging register.
// 
wire rstag_165to165_bb2_ld__u1_valid_out;
wire rstag_165to165_bb2_ld__u1_stall_in;
wire rstag_165to165_bb2_ld__u1_inputs_ready;
wire rstag_165to165_bb2_ld__u1_stall_local;
 reg rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG;
wire rstag_165to165_bb2_ld__u1_combined_valid;
 reg [31:0] rstag_165to165_bb2_ld__u1_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_165to165_bb2_ld__u1;

assign rstag_165to165_bb2_ld__u1_inputs_ready = local_bb2_ld__u1_valid_out_NO_SHIFT_REG;
assign rstag_165to165_bb2_ld__u1 = (rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG ? rstag_165to165_bb2_ld__u1_staging_reg_NO_SHIFT_REG : local_bb2_ld__u1_NO_SHIFT_REG);
assign rstag_165to165_bb2_ld__u1_combined_valid = (rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG | rstag_165to165_bb2_ld__u1_inputs_ready);
assign rstag_165to165_bb2_ld__u1_valid_out = rstag_165to165_bb2_ld__u1_combined_valid;
assign rstag_165to165_bb2_ld__u1_stall_local = rstag_165to165_bb2_ld__u1_stall_in;
assign local_bb2_ld__u1_stall_in = (|rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_165to165_bb2_ld__u1_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_165to165_bb2_ld__u1_stall_local)
		begin
			if (~(rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG))
			begin
				rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG <= rstag_165to165_bb2_ld__u1_inputs_ready;
			end
		end
		else
		begin
			rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_165to165_bb2_ld__u1_staging_valid_NO_SHIFT_REG))
		begin
			rstag_165to165_bb2_ld__u1_staging_reg_NO_SHIFT_REG <= local_bb2_ld__u1_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_ld__u2_inputs_ready;
 reg local_bb2_ld__u2_valid_out_NO_SHIFT_REG;
wire local_bb2_ld__u2_stall_in;
wire local_bb2_ld__u2_output_regs_ready;
wire local_bb2_ld__u2_fu_stall_out;
wire local_bb2_ld__u2_fu_valid_out;
wire [31:0] local_bb2_ld__u2_lsu_dataout;
 reg [31:0] local_bb2_ld__u2_NO_SHIFT_REG;
wire local_bb2_ld__u2_causedstall;

lsu_top lsu_local_bb2_ld__u2 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld__u2_fu_stall_out),
	.i_valid(local_bb2_ld__u2_inputs_ready),
	.i_address(rstag_5to5_bb2_arrayidx7_1),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rstag_5to5_bb2_cmp3_NEG_or49),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld__u2_output_regs_ready)),
	.o_valid(local_bb2_ld__u2_fu_valid_out),
	.o_readdata(local_bb2_ld__u2_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld__u2_active),
	.avm_address(avm_local_bb2_ld__u2_address),
	.avm_read(avm_local_bb2_ld__u2_read),
	.avm_readdata(avm_local_bb2_ld__u2_readdata),
	.avm_write(avm_local_bb2_ld__u2_write),
	.avm_writeack(avm_local_bb2_ld__u2_writeack),
	.avm_burstcount(avm_local_bb2_ld__u2_burstcount),
	.avm_writedata(avm_local_bb2_ld__u2_writedata),
	.avm_byteenable(avm_local_bb2_ld__u2_byteenable),
	.avm_waitrequest(avm_local_bb2_ld__u2_waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld__u2_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld__u2.AWIDTH = 30;
defparam lsu_local_bb2_ld__u2.WIDTH_BYTES = 4;
defparam lsu_local_bb2_ld__u2.MWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld__u2.WRITEDATAWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld__u2.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb2_ld__u2.READ = 1;
defparam lsu_local_bb2_ld__u2.ATOMIC = 0;
defparam lsu_local_bb2_ld__u2.WIDTH = 32;
defparam lsu_local_bb2_ld__u2.MWIDTH = 256;
defparam lsu_local_bb2_ld__u2.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld__u2.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld__u2.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld__u2.MEMORY_SIDE_MEM_LATENCY = 61;
defparam lsu_local_bb2_ld__u2.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld__u2.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld__u2.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld__u2.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld__u2.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld__u2.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld__u2.USECACHING = 1;
defparam lsu_local_bb2_ld__u2.CACHESIZE = 256;
defparam lsu_local_bb2_ld__u2.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld__u2.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld__u2.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld__u2.ADDRSPACE = 1;
defparam lsu_local_bb2_ld__u2.STYLE = "BURST-COALESCED";

assign local_bb2_ld__u2_inputs_ready = (rstag_5to5_bb2_arrayidx7_1_valid_out & rstag_5to5_bb2_cmp3_NEG_or49_valid_out_1);
assign local_bb2_ld__u2_output_regs_ready = (&(~(local_bb2_ld__u2_valid_out_NO_SHIFT_REG) | ~(local_bb2_ld__u2_stall_in)));
assign rstag_5to5_bb2_arrayidx7_1_stall_in = (local_bb2_ld__u2_fu_stall_out | ~(local_bb2_ld__u2_inputs_ready));
assign rstag_5to5_bb2_cmp3_NEG_or49_stall_in_1 = (local_bb2_ld__u2_fu_stall_out | ~(local_bb2_ld__u2_inputs_ready));
assign local_bb2_ld__u2_causedstall = (local_bb2_ld__u2_inputs_ready && (local_bb2_ld__u2_fu_stall_out && !(~(local_bb2_ld__u2_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld__u2_NO_SHIFT_REG <= 'x;
		local_bb2_ld__u2_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld__u2_output_regs_ready)
		begin
			local_bb2_ld__u2_NO_SHIFT_REG <= local_bb2_ld__u2_lsu_dataout;
			local_bb2_ld__u2_valid_out_NO_SHIFT_REG <= local_bb2_ld__u2_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld__u2_stall_in))
			begin
				local_bb2_ld__u2_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_ld__u3_inputs_ready;
 reg local_bb2_ld__u3_valid_out_NO_SHIFT_REG;
wire local_bb2_ld__u3_stall_in;
wire local_bb2_ld__u3_output_regs_ready;
wire local_bb2_ld__u3_fu_stall_out;
wire local_bb2_ld__u3_fu_valid_out;
wire [31:0] local_bb2_ld__u3_lsu_dataout;
 reg [31:0] local_bb2_ld__u3_NO_SHIFT_REG;
wire local_bb2_ld__u3_causedstall;

lsu_top lsu_local_bb2_ld__u3 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb2_ld__u3_fu_stall_out),
	.i_valid(local_bb2_ld__u3_inputs_ready),
	.i_address(rstag_5to5_bb2_arrayidx16_1),
	.i_writedata(),
	.i_cmpdata(),
	.i_predicate(rstag_5to5_bb2_cmp3_NEG_or49),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb2_ld__u3_output_regs_ready)),
	.o_valid(local_bb2_ld__u3_fu_valid_out),
	.o_readdata(local_bb2_ld__u3_lsu_dataout),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb2_ld__u3_active),
	.avm_address(avm_local_bb2_ld__u3_address),
	.avm_read(avm_local_bb2_ld__u3_read),
	.avm_readdata(avm_local_bb2_ld__u3_readdata),
	.avm_write(avm_local_bb2_ld__u3_write),
	.avm_writeack(avm_local_bb2_ld__u3_writeack),
	.avm_burstcount(avm_local_bb2_ld__u3_burstcount),
	.avm_writedata(avm_local_bb2_ld__u3_writedata),
	.avm_byteenable(avm_local_bb2_ld__u3_byteenable),
	.avm_waitrequest(avm_local_bb2_ld__u3_waitrequest),
	.avm_readdatavalid(avm_local_bb2_ld__u3_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb2_ld__u3.AWIDTH = 30;
defparam lsu_local_bb2_ld__u3.WIDTH_BYTES = 4;
defparam lsu_local_bb2_ld__u3.MWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld__u3.WRITEDATAWIDTH_BYTES = 32;
defparam lsu_local_bb2_ld__u3.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb2_ld__u3.READ = 1;
defparam lsu_local_bb2_ld__u3.ATOMIC = 0;
defparam lsu_local_bb2_ld__u3.WIDTH = 32;
defparam lsu_local_bb2_ld__u3.MWIDTH = 256;
defparam lsu_local_bb2_ld__u3.ATOMIC_WIDTH = 3;
defparam lsu_local_bb2_ld__u3.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb2_ld__u3.KERNEL_SIDE_MEM_LATENCY = 160;
defparam lsu_local_bb2_ld__u3.MEMORY_SIDE_MEM_LATENCY = 61;
defparam lsu_local_bb2_ld__u3.USE_WRITE_ACK = 0;
defparam lsu_local_bb2_ld__u3.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb2_ld__u3.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb2_ld__u3.NUMBER_BANKS = 1;
defparam lsu_local_bb2_ld__u3.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb2_ld__u3.USEINPUTFIFO = 0;
defparam lsu_local_bb2_ld__u3.USECACHING = 1;
defparam lsu_local_bb2_ld__u3.CACHESIZE = 256;
defparam lsu_local_bb2_ld__u3.USEOUTPUTFIFO = 1;
defparam lsu_local_bb2_ld__u3.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb2_ld__u3.HIGH_FMAX = 1;
defparam lsu_local_bb2_ld__u3.ADDRSPACE = 1;
defparam lsu_local_bb2_ld__u3.STYLE = "BURST-COALESCED";

assign local_bb2_ld__u3_inputs_ready = (rstag_5to5_bb2_arrayidx16_1_valid_out & rstag_5to5_bb2_cmp3_NEG_or49_valid_out_0);
assign local_bb2_ld__u3_output_regs_ready = (&(~(local_bb2_ld__u3_valid_out_NO_SHIFT_REG) | ~(local_bb2_ld__u3_stall_in)));
assign rstag_5to5_bb2_arrayidx16_1_stall_in = (local_bb2_ld__u3_fu_stall_out | ~(local_bb2_ld__u3_inputs_ready));
assign rstag_5to5_bb2_cmp3_NEG_or49_stall_in_0 = (local_bb2_ld__u3_fu_stall_out | ~(local_bb2_ld__u3_inputs_ready));
assign local_bb2_ld__u3_causedstall = (local_bb2_ld__u3_inputs_ready && (local_bb2_ld__u3_fu_stall_out && !(~(local_bb2_ld__u3_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_ld__u3_NO_SHIFT_REG <= 'x;
		local_bb2_ld__u3_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_ld__u3_output_regs_ready)
		begin
			local_bb2_ld__u3_NO_SHIFT_REG <= local_bb2_ld__u3_lsu_dataout;
			local_bb2_ld__u3_valid_out_NO_SHIFT_REG <= local_bb2_ld__u3_fu_valid_out;
		end
		else
		begin
			if (~(local_bb2_ld__u3_stall_in))
			begin
				local_bb2_ld__u3_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_c0_eni2_stall_local;
wire [351:0] local_bb2_c0_eni2;

assign local_bb2_c0_eni2[95:0] = local_bb2_c0_eni1[95:0];
assign local_bb2_c0_eni2[127:96] = rstag_165to165_bb2_ld_;
assign local_bb2_c0_eni2[351:128] = local_bb2_c0_eni1[351:128];

// This section implements a staging register.
// 
wire rstag_165to165_bb2_ld__u2_valid_out;
wire rstag_165to165_bb2_ld__u2_stall_in;
wire rstag_165to165_bb2_ld__u2_inputs_ready;
wire rstag_165to165_bb2_ld__u2_stall_local;
 reg rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG;
wire rstag_165to165_bb2_ld__u2_combined_valid;
 reg [31:0] rstag_165to165_bb2_ld__u2_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_165to165_bb2_ld__u2;

assign rstag_165to165_bb2_ld__u2_inputs_ready = local_bb2_ld__u2_valid_out_NO_SHIFT_REG;
assign rstag_165to165_bb2_ld__u2 = (rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG ? rstag_165to165_bb2_ld__u2_staging_reg_NO_SHIFT_REG : local_bb2_ld__u2_NO_SHIFT_REG);
assign rstag_165to165_bb2_ld__u2_combined_valid = (rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG | rstag_165to165_bb2_ld__u2_inputs_ready);
assign rstag_165to165_bb2_ld__u2_valid_out = rstag_165to165_bb2_ld__u2_combined_valid;
assign rstag_165to165_bb2_ld__u2_stall_local = rstag_165to165_bb2_ld__u2_stall_in;
assign local_bb2_ld__u2_stall_in = (|rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_165to165_bb2_ld__u2_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_165to165_bb2_ld__u2_stall_local)
		begin
			if (~(rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG))
			begin
				rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG <= rstag_165to165_bb2_ld__u2_inputs_ready;
			end
		end
		else
		begin
			rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_165to165_bb2_ld__u2_staging_valid_NO_SHIFT_REG))
		begin
			rstag_165to165_bb2_ld__u2_staging_reg_NO_SHIFT_REG <= local_bb2_ld__u2_NO_SHIFT_REG;
		end
	end
end


// This section implements a staging register.
// 
wire rstag_165to165_bb2_ld__u3_valid_out;
wire rstag_165to165_bb2_ld__u3_stall_in;
wire rstag_165to165_bb2_ld__u3_inputs_ready;
wire rstag_165to165_bb2_ld__u3_stall_local;
 reg rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG;
wire rstag_165to165_bb2_ld__u3_combined_valid;
 reg [31:0] rstag_165to165_bb2_ld__u3_staging_reg_NO_SHIFT_REG;
wire [31:0] rstag_165to165_bb2_ld__u3;

assign rstag_165to165_bb2_ld__u3_inputs_ready = local_bb2_ld__u3_valid_out_NO_SHIFT_REG;
assign rstag_165to165_bb2_ld__u3 = (rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG ? rstag_165to165_bb2_ld__u3_staging_reg_NO_SHIFT_REG : local_bb2_ld__u3_NO_SHIFT_REG);
assign rstag_165to165_bb2_ld__u3_combined_valid = (rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG | rstag_165to165_bb2_ld__u3_inputs_ready);
assign rstag_165to165_bb2_ld__u3_valid_out = rstag_165to165_bb2_ld__u3_combined_valid;
assign rstag_165to165_bb2_ld__u3_stall_local = rstag_165to165_bb2_ld__u3_stall_in;
assign local_bb2_ld__u3_stall_in = (|rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_165to165_bb2_ld__u3_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_165to165_bb2_ld__u3_stall_local)
		begin
			if (~(rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG))
			begin
				rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG <= rstag_165to165_bb2_ld__u3_inputs_ready;
			end
		end
		else
		begin
			rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_165to165_bb2_ld__u3_staging_valid_NO_SHIFT_REG))
		begin
			rstag_165to165_bb2_ld__u3_staging_reg_NO_SHIFT_REG <= local_bb2_ld__u3_NO_SHIFT_REG;
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_c0_eni3_stall_local;
wire [351:0] local_bb2_c0_eni3;

assign local_bb2_c0_eni3[127:0] = local_bb2_c0_eni2[127:0];
assign local_bb2_c0_eni3[191:128] = rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_NO_SHIFT_REG;
assign local_bb2_c0_eni3[351:192] = local_bb2_c0_eni2[351:192];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_eni4_stall_local;
wire [351:0] local_bb2_c0_eni4;

assign local_bb2_c0_eni4[191:0] = local_bb2_c0_eni3[191:0];
assign local_bb2_c0_eni4[223:192] = rstag_165to165_bb2_ld__u1;
assign local_bb2_c0_eni4[351:224] = local_bb2_c0_eni3[351:224];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_eni5_stall_local;
wire [351:0] local_bb2_c0_eni5;

assign local_bb2_c0_eni5[223:0] = local_bb2_c0_eni4[223:0];
assign local_bb2_c0_eni5[255:224] = rnode_164to165_tmpr_05_0_NO_SHIFT_REG;
assign local_bb2_c0_eni5[351:256] = local_bb2_c0_eni4[351:256];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_eni6_stall_local;
wire [351:0] local_bb2_c0_eni6;

assign local_bb2_c0_eni6[255:0] = local_bb2_c0_eni5[255:0];
assign local_bb2_c0_eni6[287:256] = rnode_164to165_tmpi_06_0_NO_SHIFT_REG;
assign local_bb2_c0_eni6[351:288] = local_bb2_c0_eni5[351:288];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_eni7_stall_local;
wire [351:0] local_bb2_c0_eni7;

assign local_bb2_c0_eni7[287:0] = local_bb2_c0_eni6[287:0];
assign local_bb2_c0_eni7[319:288] = rstag_165to165_bb2_ld__u2;
assign local_bb2_c0_eni7[351:320] = local_bb2_c0_eni6[351:320];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_eni8_valid_out;
wire local_bb2_c0_eni8_stall_in;
wire local_bb2_c0_eni8_inputs_ready;
wire local_bb2_c0_eni8_stall_local;
wire [351:0] local_bb2_c0_eni8;

assign local_bb2_c0_eni8_inputs_ready = (rnode_164to165_tmpr_05_0_valid_out_NO_SHIFT_REG & rnode_164to165_tmpi_06_0_valid_out_NO_SHIFT_REG & rstag_165to165_bb2_ld__u2_valid_out & rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_valid_out_NO_SHIFT_REG & rstag_165to165_bb2_ld__valid_out & rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_valid_out_NO_SHIFT_REG & rstag_165to165_bb2_ld__u1_valid_out & rstag_165to165_bb2_ld__u3_valid_out);
assign local_bb2_c0_eni8[319:0] = local_bb2_c0_eni7[319:0];
assign local_bb2_c0_eni8[351:320] = rstag_165to165_bb2_ld__u3;
assign local_bb2_c0_eni8_valid_out = local_bb2_c0_eni8_inputs_ready;
assign local_bb2_c0_eni8_stall_local = local_bb2_c0_eni8_stall_in;
assign rnode_164to165_tmpr_05_0_stall_in_NO_SHIFT_REG = (local_bb2_c0_eni8_stall_local | ~(local_bb2_c0_eni8_inputs_ready));
assign rnode_164to165_tmpi_06_0_stall_in_NO_SHIFT_REG = (local_bb2_c0_eni8_stall_local | ~(local_bb2_c0_eni8_inputs_ready));
assign rstag_165to165_bb2_ld__u2_stall_in = (local_bb2_c0_eni8_stall_local | ~(local_bb2_c0_eni8_inputs_ready));
assign rnode_165to165_bb2_ld_memcoalesce_m1r_load_0_0_stall_in_NO_SHIFT_REG = (local_bb2_c0_eni8_stall_local | ~(local_bb2_c0_eni8_inputs_ready));
assign rstag_165to165_bb2_ld__stall_in = (local_bb2_c0_eni8_stall_local | ~(local_bb2_c0_eni8_inputs_ready));
assign rnode_165to165_bb2_ld_memcoalesce_m1i_load_0_0_stall_in_NO_SHIFT_REG = (local_bb2_c0_eni8_stall_local | ~(local_bb2_c0_eni8_inputs_ready));
assign rstag_165to165_bb2_ld__u1_stall_in = (local_bb2_c0_eni8_stall_local | ~(local_bb2_c0_eni8_inputs_ready));
assign rstag_165to165_bb2_ld__u3_stall_in = (local_bb2_c0_eni8_stall_local | ~(local_bb2_c0_eni8_inputs_ready));

// This section implements a registered operation.
// 
wire local_bb2_c0_enter_c0_eni8_inputs_ready;
 reg local_bb2_c0_enter_c0_eni8_valid_out_0_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_stall_in_0;
 reg local_bb2_c0_enter_c0_eni8_valid_out_1_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_stall_in_1;
 reg local_bb2_c0_enter_c0_eni8_valid_out_2_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_stall_in_2;
 reg local_bb2_c0_enter_c0_eni8_valid_out_3_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_stall_in_3;
 reg local_bb2_c0_enter_c0_eni8_valid_out_4_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_stall_in_4;
 reg local_bb2_c0_enter_c0_eni8_valid_out_5_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_stall_in_5;
 reg local_bb2_c0_enter_c0_eni8_valid_out_6_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_stall_in_6;
 reg local_bb2_c0_enter_c0_eni8_valid_out_7_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_stall_in_7;
wire local_bb2_c0_enter_c0_eni8_output_regs_ready;
 reg [351:0] local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG;
wire local_bb2_c0_enter_c0_eni8_input_accepted;
wire local_bb2_c0_exit_c0_exi4_entry_stall;
wire local_bb2_c0_exit_c0_exi4_output_regs_ready;
wire [26:0] local_bb2_c0_exit_c0_exi4_valid_bits;
wire local_bb2_c0_exit_c0_exi4_phases;
wire local_bb2_c0_enter_c0_eni8_inc_pipelined_thread;
wire local_bb2_c0_enter_c0_eni8_dec_pipelined_thread;
wire local_bb2_c0_enter_c0_eni8_causedstall;

assign local_bb2_c0_enter_c0_eni8_inputs_ready = local_bb2_c0_eni8_valid_out;
assign local_bb2_c0_enter_c0_eni8_output_regs_ready = 1'b1;
assign local_bb2_c0_enter_c0_eni8_input_accepted = (local_bb2_c0_enter_c0_eni8_inputs_ready && !(local_bb2_c0_exit_c0_exi4_entry_stall));
assign local_bb2_c0_enter_c0_eni8_inc_pipelined_thread = 1'b1;
assign local_bb2_c0_enter_c0_eni8_dec_pipelined_thread = ~(1'b0);
assign local_bb2_c0_eni8_stall_in = ((~(local_bb2_c0_enter_c0_eni8_inputs_ready) | local_bb2_c0_exit_c0_exi4_entry_stall) | ~(1'b1));
assign local_bb2_c0_enter_c0_eni8_causedstall = (1'b1 && ((~(local_bb2_c0_enter_c0_eni8_inputs_ready) | local_bb2_c0_exit_c0_exi4_entry_stall) && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG <= 'x;
		local_bb2_c0_enter_c0_eni8_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_enter_c0_eni8_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_enter_c0_eni8_valid_out_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_enter_c0_eni8_valid_out_3_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_enter_c0_eni8_valid_out_4_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_enter_c0_eni8_valid_out_5_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_enter_c0_eni8_valid_out_6_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_enter_c0_eni8_valid_out_7_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_c0_enter_c0_eni8_output_regs_ready)
		begin
			local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG <= local_bb2_c0_eni8;
			local_bb2_c0_enter_c0_eni8_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_c0_enter_c0_eni8_valid_out_1_NO_SHIFT_REG <= 1'b1;
			local_bb2_c0_enter_c0_eni8_valid_out_2_NO_SHIFT_REG <= 1'b1;
			local_bb2_c0_enter_c0_eni8_valid_out_3_NO_SHIFT_REG <= 1'b1;
			local_bb2_c0_enter_c0_eni8_valid_out_4_NO_SHIFT_REG <= 1'b1;
			local_bb2_c0_enter_c0_eni8_valid_out_5_NO_SHIFT_REG <= 1'b1;
			local_bb2_c0_enter_c0_eni8_valid_out_6_NO_SHIFT_REG <= 1'b1;
			local_bb2_c0_enter_c0_eni8_valid_out_7_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_c0_enter_c0_eni8_stall_in_0))
			begin
				local_bb2_c0_enter_c0_eni8_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_enter_c0_eni8_stall_in_1))
			begin
				local_bb2_c0_enter_c0_eni8_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_enter_c0_eni8_stall_in_2))
			begin
				local_bb2_c0_enter_c0_eni8_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_enter_c0_eni8_stall_in_3))
			begin
				local_bb2_c0_enter_c0_eni8_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_enter_c0_eni8_stall_in_4))
			begin
				local_bb2_c0_enter_c0_eni8_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_enter_c0_eni8_stall_in_5))
			begin
				local_bb2_c0_enter_c0_eni8_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_enter_c0_eni8_stall_in_6))
			begin
				local_bb2_c0_enter_c0_eni8_valid_out_6_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_enter_c0_eni8_stall_in_7))
			begin
				local_bb2_c0_enter_c0_eni8_valid_out_7_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_c0_ene1_stall_local;
wire [63:0] local_bb2_c0_ene1;

assign local_bb2_c0_ene1 = local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG[95:32];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_ene2_stall_local;
wire [31:0] local_bb2_c0_ene2;

assign local_bb2_c0_ene2 = local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG[127:96];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_ene3_stall_local;
wire [63:0] local_bb2_c0_ene3;

assign local_bb2_c0_ene3 = local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG[191:128];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_ene4_stall_local;
wire [31:0] local_bb2_c0_ene4;

assign local_bb2_c0_ene4 = local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG[223:192];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_ene5_valid_out;
wire local_bb2_c0_ene5_stall_in;
wire local_bb2_c0_ene5_inputs_ready;
wire local_bb2_c0_ene5_stall_local;
wire [31:0] local_bb2_c0_ene5;

assign local_bb2_c0_ene5_inputs_ready = local_bb2_c0_enter_c0_eni8_valid_out_4_NO_SHIFT_REG;
assign local_bb2_c0_ene5 = local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG[255:224];
assign local_bb2_c0_ene5_valid_out = 1'b1;
assign local_bb2_c0_enter_c0_eni8_stall_in_4 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_c0_ene6_valid_out;
wire local_bb2_c0_ene6_stall_in;
wire local_bb2_c0_ene6_inputs_ready;
wire local_bb2_c0_ene6_stall_local;
wire [31:0] local_bb2_c0_ene6;

assign local_bb2_c0_ene6_inputs_ready = local_bb2_c0_enter_c0_eni8_valid_out_5_NO_SHIFT_REG;
assign local_bb2_c0_ene6 = local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG[287:256];
assign local_bb2_c0_ene6_valid_out = 1'b1;
assign local_bb2_c0_enter_c0_eni8_stall_in_5 = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_c0_ene7_stall_local;
wire [31:0] local_bb2_c0_ene7;

assign local_bb2_c0_ene7 = local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG[319:288];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_ene8_stall_local;
wire [31:0] local_bb2_c0_ene8;

assign local_bb2_c0_ene8 = local_bb2_c0_enter_c0_eni8_NO_SHIFT_REG[351:320];

// This section implements an unregistered operation.
// 
wire local_bb2_memcoalesce_m1r_extrValue_0_stall_local;
wire [31:0] local_bb2_memcoalesce_m1r_extrValue_0;

assign local_bb2_memcoalesce_m1r_extrValue_0 = local_bb2_c0_ene1[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_memcoalesce_m1r_extrValue_1_stall_local;
wire [31:0] local_bb2_memcoalesce_m1r_extrValue_1;

assign local_bb2_memcoalesce_m1r_extrValue_1 = local_bb2_c0_ene1[63:32];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u4_stall_local;
wire [31:0] local_bb2_var__u4;

assign local_bb2_var__u4 = local_bb2_c0_ene2;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u5_stall_local;
wire [31:0] local_bb2_var__u5;

assign local_bb2_var__u5 = local_bb2_c0_ene2;

// This section implements an unregistered operation.
// 
wire local_bb2_memcoalesce_m1i_extrValue_0_stall_local;
wire [31:0] local_bb2_memcoalesce_m1i_extrValue_0;

assign local_bb2_memcoalesce_m1i_extrValue_0 = local_bb2_c0_ene3[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_memcoalesce_m1i_extrValue_1_stall_local;
wire [31:0] local_bb2_memcoalesce_m1i_extrValue_1;

assign local_bb2_memcoalesce_m1i_extrValue_1 = local_bb2_c0_ene3[63:32];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u6_stall_local;
wire [31:0] local_bb2_var__u6;

assign local_bb2_var__u6 = local_bb2_c0_ene4;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u7_stall_local;
wire [31:0] local_bb2_var__u7;

assign local_bb2_var__u7 = local_bb2_c0_ene4;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene5_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_c0_ene5_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene5_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene5_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene5_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_c0_ene5_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_c0_ene5_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_c0_ene5_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_c0_ene5_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_c0_ene5_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_c0_ene5),
	.data_out(rnode_166to167_bb2_c0_ene5_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_c0_ene5_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_c0_ene5_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_c0_ene5_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_c0_ene5_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_c0_ene5_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_c0_ene5_stall_in = 1'b0;
assign rnode_166to167_bb2_c0_ene5_0_NO_SHIFT_REG = rnode_166to167_bb2_c0_ene5_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_c0_ene5_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene6_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_c0_ene6_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene6_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene6_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_c0_ene6_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_c0_ene6_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_c0_ene6_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_c0_ene6_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_c0_ene6_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_c0_ene6_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_c0_ene6),
	.data_out(rnode_166to167_bb2_c0_ene6_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_c0_ene6_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_c0_ene6_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_c0_ene6_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_c0_ene6_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_c0_ene6_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_c0_ene6_stall_in = 1'b0;
assign rnode_166to167_bb2_c0_ene6_0_NO_SHIFT_REG = rnode_166to167_bb2_c0_ene6_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_c0_ene6_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u8_stall_local;
wire [31:0] local_bb2_var__u8;

assign local_bb2_var__u8 = local_bb2_c0_ene7;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u9_stall_local;
wire [31:0] local_bb2_var__u9;

assign local_bb2_var__u9 = local_bb2_c0_ene7;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u10_stall_local;
wire [31:0] local_bb2_var__u10;

assign local_bb2_var__u10 = local_bb2_c0_ene8;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u11_stall_local;
wire [31:0] local_bb2_var__u11;

assign local_bb2_var__u11 = local_bb2_c0_ene8;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u12_stall_local;
wire [31:0] local_bb2_var__u12;

assign local_bb2_var__u12 = local_bb2_memcoalesce_m1r_extrValue_0;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u13_stall_local;
wire [31:0] local_bb2_var__u13;

assign local_bb2_var__u13 = local_bb2_memcoalesce_m1r_extrValue_0;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u14_stall_local;
wire [31:0] local_bb2_var__u14;

assign local_bb2_var__u14 = local_bb2_memcoalesce_m1r_extrValue_1;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u15_stall_local;
wire [31:0] local_bb2_var__u15;

assign local_bb2_var__u15 = local_bb2_memcoalesce_m1r_extrValue_1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr2_i_stall_local;
wire [31:0] local_bb2_shr2_i;

assign local_bb2_shr2_i = (local_bb2_var__u4 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and6_i_stall_local;
wire [31:0] local_bb2_and6_i;

assign local_bb2_and6_i = (local_bb2_var__u4 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr2_i1276_stall_local;
wire [31:0] local_bb2_shr2_i1276;

assign local_bb2_shr2_i1276 = (local_bb2_var__u5 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and6_i1281_stall_local;
wire [31:0] local_bb2_and6_i1281;

assign local_bb2_and6_i1281 = (local_bb2_var__u5 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u16_stall_local;
wire [31:0] local_bb2_var__u16;

assign local_bb2_var__u16 = local_bb2_memcoalesce_m1i_extrValue_0;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u17_stall_local;
wire [31:0] local_bb2_var__u17;

assign local_bb2_var__u17 = local_bb2_memcoalesce_m1i_extrValue_0;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u18_stall_local;
wire [31:0] local_bb2_var__u18;

assign local_bb2_var__u18 = local_bb2_memcoalesce_m1i_extrValue_1;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u19_stall_local;
wire [31:0] local_bb2_var__u19;

assign local_bb2_var__u19 = local_bb2_memcoalesce_m1i_extrValue_1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr2_i1825_stall_local;
wire [31:0] local_bb2_shr2_i1825;

assign local_bb2_shr2_i1825 = (local_bb2_var__u6 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and6_i1830_stall_local;
wire [31:0] local_bb2_and6_i1830;

assign local_bb2_and6_i1830 = (local_bb2_var__u6 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr2_i1368_stall_local;
wire [31:0] local_bb2_shr2_i1368;

assign local_bb2_shr2_i1368 = (local_bb2_var__u7 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and6_i1373_stall_local;
wire [31:0] local_bb2_and6_i1373;

assign local_bb2_and6_i1373 = (local_bb2_var__u7 & 32'h7FFFFF);

// Register node:
//  * latency = 10
//  * capacity = 10
 logic rnode_167to177_bb2_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to177_bb2_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene5_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to177_bb2_c0_ene5_0_reg_177_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene5_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene5_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene5_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_167to177_bb2_c0_ene5_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to177_bb2_c0_ene5_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to177_bb2_c0_ene5_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_167to177_bb2_c0_ene5_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_167to177_bb2_c0_ene5_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_167to177_bb2_c0_ene5_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_167to177_bb2_c0_ene5_0_reg_177_fifo.DEPTH = 10;
defparam rnode_167to177_bb2_c0_ene5_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_167to177_bb2_c0_ene5_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to177_bb2_c0_ene5_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_167to177_bb2_c0_ene5_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to177_bb2_c0_ene5_0_NO_SHIFT_REG = rnode_167to177_bb2_c0_ene5_0_reg_177_NO_SHIFT_REG;
assign rnode_167to177_bb2_c0_ene5_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_167to177_bb2_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 10
//  * capacity = 10
 logic rnode_167to177_bb2_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to177_bb2_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene6_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to177_bb2_c0_ene6_0_reg_177_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene6_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene6_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_167to177_bb2_c0_ene6_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_167to177_bb2_c0_ene6_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to177_bb2_c0_ene6_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to177_bb2_c0_ene6_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_167to177_bb2_c0_ene6_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_167to177_bb2_c0_ene6_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_c0_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_167to177_bb2_c0_ene6_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_167to177_bb2_c0_ene6_0_reg_177_fifo.DEPTH = 10;
defparam rnode_167to177_bb2_c0_ene6_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_167to177_bb2_c0_ene6_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to177_bb2_c0_ene6_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_167to177_bb2_c0_ene6_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to177_bb2_c0_ene6_0_NO_SHIFT_REG = rnode_167to177_bb2_c0_ene6_0_reg_177_NO_SHIFT_REG;
assign rnode_167to177_bb2_c0_ene6_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_167to177_bb2_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr2_i820_stall_local;
wire [31:0] local_bb2_shr2_i820;

assign local_bb2_shr2_i820 = (local_bb2_var__u8 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and6_i825_stall_local;
wire [31:0] local_bb2_and6_i825;

assign local_bb2_and6_i825 = (local_bb2_var__u8 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr2_i264_stall_local;
wire [31:0] local_bb2_shr2_i264;

assign local_bb2_shr2_i264 = (local_bb2_var__u9 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and6_i269_stall_local;
wire [31:0] local_bb2_and6_i269;

assign local_bb2_and6_i269 = (local_bb2_var__u9 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr2_i728_stall_local;
wire [31:0] local_bb2_shr2_i728;

assign local_bb2_shr2_i728 = (local_bb2_var__u10 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and6_i733_stall_local;
wire [31:0] local_bb2_and6_i733;

assign local_bb2_and6_i733 = (local_bb2_var__u10 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr2_i356_stall_local;
wire [31:0] local_bb2_shr2_i356;

assign local_bb2_shr2_i356 = (local_bb2_var__u11 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and6_i361_stall_local;
wire [31:0] local_bb2_and6_i361;

assign local_bb2_and6_i361 = (local_bb2_var__u11 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_stall_local;
wire [31:0] local_bb2_shr_i;

assign local_bb2_shr_i = (local_bb2_var__u12 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i_stall_local;
wire [31:0] local_bb2_xor_i;

assign local_bb2_xor_i = (local_bb2_var__u4 ^ local_bb2_var__u12);

// This section implements an unregistered operation.
// 
wire local_bb2_and5_i_stall_local;
wire [31:0] local_bb2_and5_i;

assign local_bb2_and5_i = (local_bb2_var__u12 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i1366_stall_local;
wire [31:0] local_bb2_shr_i1366;

assign local_bb2_shr_i1366 = (local_bb2_var__u13 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i1370_stall_local;
wire [31:0] local_bb2_xor_i1370;

assign local_bb2_xor_i1370 = (local_bb2_var__u7 ^ local_bb2_var__u13);

// This section implements an unregistered operation.
// 
wire local_bb2_and5_i1372_stall_local;
wire [31:0] local_bb2_and5_i1372;

assign local_bb2_and5_i1372 = (local_bb2_var__u13 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i818_stall_local;
wire [31:0] local_bb2_shr_i818;

assign local_bb2_shr_i818 = (local_bb2_var__u14 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i822_stall_local;
wire [31:0] local_bb2_xor_i822;

assign local_bb2_xor_i822 = (local_bb2_var__u8 ^ local_bb2_var__u14);

// This section implements an unregistered operation.
// 
wire local_bb2_and5_i824_stall_local;
wire [31:0] local_bb2_and5_i824;

assign local_bb2_and5_i824 = (local_bb2_var__u14 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i354_stall_local;
wire [31:0] local_bb2_shr_i354;

assign local_bb2_shr_i354 = (local_bb2_var__u15 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i358_stall_local;
wire [31:0] local_bb2_xor_i358;

assign local_bb2_xor_i358 = (local_bb2_var__u11 ^ local_bb2_var__u15);

// This section implements an unregistered operation.
// 
wire local_bb2_and5_i360_stall_local;
wire [31:0] local_bb2_and5_i360;

assign local_bb2_and5_i360 = (local_bb2_var__u15 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and3_i_stall_local;
wire [31:0] local_bb2_and3_i;

assign local_bb2_and3_i = (local_bb2_shr2_i & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_i_stall_local;
wire local_bb2_lnot17_i;

assign local_bb2_lnot17_i = (local_bb2_and6_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or47_i_stall_local;
wire [31:0] local_bb2_or47_i;

assign local_bb2_or47_i = (local_bb2_and6_i | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and3_i1277_stall_local;
wire [31:0] local_bb2_and3_i1277;

assign local_bb2_and3_i1277 = (local_bb2_shr2_i1276 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_i1287_stall_local;
wire local_bb2_lnot17_i1287;

assign local_bb2_lnot17_i1287 = (local_bb2_and6_i1281 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or47_i1309_stall_local;
wire [31:0] local_bb2_or47_i1309;

assign local_bb2_or47_i1309 = (local_bb2_and6_i1281 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i1823_stall_local;
wire [31:0] local_bb2_shr_i1823;

assign local_bb2_shr_i1823 = (local_bb2_var__u16 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i1827_stall_local;
wire [31:0] local_bb2_xor_i1827;

assign local_bb2_xor_i1827 = (local_bb2_var__u6 ^ local_bb2_var__u16);

// This section implements an unregistered operation.
// 
wire local_bb2_and5_i1829_stall_local;
wire [31:0] local_bb2_and5_i1829;

assign local_bb2_and5_i1829 = (local_bb2_var__u16 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i1274_stall_local;
wire [31:0] local_bb2_shr_i1274;

assign local_bb2_shr_i1274 = (local_bb2_var__u17 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i1278_stall_local;
wire [31:0] local_bb2_xor_i1278;

assign local_bb2_xor_i1278 = (local_bb2_var__u5 ^ local_bb2_var__u17);

// This section implements an unregistered operation.
// 
wire local_bb2_and5_i1280_stall_local;
wire [31:0] local_bb2_and5_i1280;

assign local_bb2_and5_i1280 = (local_bb2_var__u17 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i726_stall_local;
wire [31:0] local_bb2_shr_i726;

assign local_bb2_shr_i726 = (local_bb2_var__u18 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i730_stall_local;
wire [31:0] local_bb2_xor_i730;

assign local_bb2_xor_i730 = (local_bb2_var__u10 ^ local_bb2_var__u18);

// This section implements an unregistered operation.
// 
wire local_bb2_and5_i732_stall_local;
wire [31:0] local_bb2_and5_i732;

assign local_bb2_and5_i732 = (local_bb2_var__u18 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i262_stall_local;
wire [31:0] local_bb2_shr_i262;

assign local_bb2_shr_i262 = (local_bb2_var__u19 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i266_stall_local;
wire [31:0] local_bb2_xor_i266;

assign local_bb2_xor_i266 = (local_bb2_var__u9 ^ local_bb2_var__u19);

// This section implements an unregistered operation.
// 
wire local_bb2_and5_i268_stall_local;
wire [31:0] local_bb2_and5_i268;

assign local_bb2_and5_i268 = (local_bb2_var__u19 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and3_i1826_stall_local;
wire [31:0] local_bb2_and3_i1826;

assign local_bb2_and3_i1826 = (local_bb2_shr2_i1825 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_i1836_stall_local;
wire local_bb2_lnot17_i1836;

assign local_bb2_lnot17_i1836 = (local_bb2_and6_i1830 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or47_i1858_stall_local;
wire [31:0] local_bb2_or47_i1858;

assign local_bb2_or47_i1858 = (local_bb2_and6_i1830 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and3_i1369_stall_local;
wire [31:0] local_bb2_and3_i1369;

assign local_bb2_and3_i1369 = (local_bb2_shr2_i1368 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_i1379_stall_local;
wire local_bb2_lnot17_i1379;

assign local_bb2_lnot17_i1379 = (local_bb2_and6_i1373 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or47_i1401_stall_local;
wire [31:0] local_bb2_or47_i1401;

assign local_bb2_or47_i1401 = (local_bb2_and6_i1373 | 32'h800000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb2_c0_ene5_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene5_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_c0_ene5_0_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene5_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_c0_ene5_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene5_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene5_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene5_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb2_c0_ene5_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb2_c0_ene5_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb2_c0_ene5_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb2_c0_ene5_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb2_c0_ene5_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(rnode_167to177_bb2_c0_ene5_0_NO_SHIFT_REG),
	.data_out(rnode_177to178_bb2_c0_ene5_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb2_c0_ene5_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb2_c0_ene5_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb2_c0_ene5_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb2_c0_ene5_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb2_c0_ene5_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to177_bb2_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_c0_ene5_0_NO_SHIFT_REG = rnode_177to178_bb2_c0_ene5_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_c0_ene5_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_c0_ene5_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb2_c0_ene6_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene6_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_c0_ene6_0_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene6_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_c0_ene6_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene6_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene6_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_c0_ene6_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb2_c0_ene6_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb2_c0_ene6_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb2_c0_ene6_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb2_c0_ene6_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb2_c0_ene6_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(rnode_167to177_bb2_c0_ene6_0_NO_SHIFT_REG),
	.data_out(rnode_177to178_bb2_c0_ene6_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb2_c0_ene6_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb2_c0_ene6_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb2_c0_ene6_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb2_c0_ene6_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb2_c0_ene6_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to177_bb2_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_c0_ene6_0_NO_SHIFT_REG = rnode_177to178_bb2_c0_ene6_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_c0_ene6_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_c0_ene6_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and3_i821_stall_local;
wire [31:0] local_bb2_and3_i821;

assign local_bb2_and3_i821 = (local_bb2_shr2_i820 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_i831_stall_local;
wire local_bb2_lnot17_i831;

assign local_bb2_lnot17_i831 = (local_bb2_and6_i825 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or47_i853_stall_local;
wire [31:0] local_bb2_or47_i853;

assign local_bb2_or47_i853 = (local_bb2_and6_i825 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and3_i265_stall_local;
wire [31:0] local_bb2_and3_i265;

assign local_bb2_and3_i265 = (local_bb2_shr2_i264 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_i275_stall_local;
wire local_bb2_lnot17_i275;

assign local_bb2_lnot17_i275 = (local_bb2_and6_i269 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or47_i297_stall_local;
wire [31:0] local_bb2_or47_i297;

assign local_bb2_or47_i297 = (local_bb2_and6_i269 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and3_i729_stall_local;
wire [31:0] local_bb2_and3_i729;

assign local_bb2_and3_i729 = (local_bb2_shr2_i728 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_i739_stall_local;
wire local_bb2_lnot17_i739;

assign local_bb2_lnot17_i739 = (local_bb2_and6_i733 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or47_i761_stall_local;
wire [31:0] local_bb2_or47_i761;

assign local_bb2_or47_i761 = (local_bb2_and6_i733 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and3_i357_stall_local;
wire [31:0] local_bb2_and3_i357;

assign local_bb2_and3_i357 = (local_bb2_shr2_i356 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_i367_stall_local;
wire local_bb2_lnot17_i367;

assign local_bb2_lnot17_i367 = (local_bb2_and6_i361 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or47_i389_stall_local;
wire [31:0] local_bb2_or47_i389;

assign local_bb2_or47_i389 = (local_bb2_and6_i361 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_stall_local;
wire [31:0] local_bb2_and_i;

assign local_bb2_and_i = (local_bb2_shr_i & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_i_stall_local;
wire local_bb2_lnot14_i;

assign local_bb2_lnot14_i = (local_bb2_and5_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_stall_local;
wire [31:0] local_bb2_or_i;

assign local_bb2_or_i = (local_bb2_and5_i | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i1367_stall_local;
wire [31:0] local_bb2_and_i1367;

assign local_bb2_and_i1367 = (local_bb2_shr_i1366 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_i1378_stall_local;
wire local_bb2_lnot14_i1378;

assign local_bb2_lnot14_i1378 = (local_bb2_and5_i1372 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i1400_stall_local;
wire [31:0] local_bb2_or_i1400;

assign local_bb2_or_i1400 = (local_bb2_and5_i1372 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i819_stall_local;
wire [31:0] local_bb2_and_i819;

assign local_bb2_and_i819 = (local_bb2_shr_i818 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_i830_stall_local;
wire local_bb2_lnot14_i830;

assign local_bb2_lnot14_i830 = (local_bb2_and5_i824 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i852_stall_local;
wire [31:0] local_bb2_or_i852;

assign local_bb2_or_i852 = (local_bb2_and5_i824 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i355_stall_local;
wire [31:0] local_bb2_and_i355;

assign local_bb2_and_i355 = (local_bb2_shr_i354 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_i366_stall_local;
wire local_bb2_lnot14_i366;

assign local_bb2_lnot14_i366 = (local_bb2_and5_i360 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i388_stall_local;
wire [31:0] local_bb2_or_i388;

assign local_bb2_or_i388 = (local_bb2_and5_i360 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot8_i_stall_local;
wire local_bb2_lnot8_i;

assign local_bb2_lnot8_i = (local_bb2_and3_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_i_stall_local;
wire local_bb2_cmp11_i;

assign local_bb2_cmp11_i = (local_bb2_and3_i == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u20_stall_local;
wire [31:0] local_bb2_var__u20;

assign local_bb2_var__u20 = (local_bb2_and3_i | local_bb2_and6_i);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_not_i_stall_local;
wire local_bb2_lnot17_not_i;

assign local_bb2_lnot17_not_i = (local_bb2_lnot17_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv1_i_i_stall_local;
wire [63:0] local_bb2_conv1_i_i;

assign local_bb2_conv1_i_i[63:32] = 32'h0;
assign local_bb2_conv1_i_i[31:0] = local_bb2_or47_i;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot8_i1283_stall_local;
wire local_bb2_lnot8_i1283;

assign local_bb2_lnot8_i1283 = (local_bb2_and3_i1277 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_i1285_stall_local;
wire local_bb2_cmp11_i1285;

assign local_bb2_cmp11_i1285 = (local_bb2_and3_i1277 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u21_stall_local;
wire [31:0] local_bb2_var__u21;

assign local_bb2_var__u21 = (local_bb2_and3_i1277 | local_bb2_and6_i1281);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_not_i1291_stall_local;
wire local_bb2_lnot17_not_i1291;

assign local_bb2_lnot17_not_i1291 = (local_bb2_lnot17_i1287 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv1_i_i1311_stall_local;
wire [63:0] local_bb2_conv1_i_i1311;

assign local_bb2_conv1_i_i1311[63:32] = 32'h0;
assign local_bb2_conv1_i_i1311[31:0] = local_bb2_or47_i1309;

// This section implements an unregistered operation.
// 
wire local_bb2_and_i1824_stall_local;
wire [31:0] local_bb2_and_i1824;

assign local_bb2_and_i1824 = (local_bb2_shr_i1823 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_i1835_stall_local;
wire local_bb2_lnot14_i1835;

assign local_bb2_lnot14_i1835 = (local_bb2_and5_i1829 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i1857_stall_local;
wire [31:0] local_bb2_or_i1857;

assign local_bb2_or_i1857 = (local_bb2_and5_i1829 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i1275_stall_local;
wire [31:0] local_bb2_and_i1275;

assign local_bb2_and_i1275 = (local_bb2_shr_i1274 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_i1286_stall_local;
wire local_bb2_lnot14_i1286;

assign local_bb2_lnot14_i1286 = (local_bb2_and5_i1280 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i1308_stall_local;
wire [31:0] local_bb2_or_i1308;

assign local_bb2_or_i1308 = (local_bb2_and5_i1280 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i727_stall_local;
wire [31:0] local_bb2_and_i727;

assign local_bb2_and_i727 = (local_bb2_shr_i726 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_i738_stall_local;
wire local_bb2_lnot14_i738;

assign local_bb2_lnot14_i738 = (local_bb2_and5_i732 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i760_stall_local;
wire [31:0] local_bb2_or_i760;

assign local_bb2_or_i760 = (local_bb2_and5_i732 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i263_stall_local;
wire [31:0] local_bb2_and_i263;

assign local_bb2_and_i263 = (local_bb2_shr_i262 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_i274_stall_local;
wire local_bb2_lnot14_i274;

assign local_bb2_lnot14_i274 = (local_bb2_and5_i268 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i296_stall_local;
wire [31:0] local_bb2_or_i296;

assign local_bb2_or_i296 = (local_bb2_and5_i268 | 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot8_i1832_stall_local;
wire local_bb2_lnot8_i1832;

assign local_bb2_lnot8_i1832 = (local_bb2_and3_i1826 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_i1834_stall_local;
wire local_bb2_cmp11_i1834;

assign local_bb2_cmp11_i1834 = (local_bb2_and3_i1826 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u22_stall_local;
wire [31:0] local_bb2_var__u22;

assign local_bb2_var__u22 = (local_bb2_and3_i1826 | local_bb2_and6_i1830);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_not_i1840_stall_local;
wire local_bb2_lnot17_not_i1840;

assign local_bb2_lnot17_not_i1840 = (local_bb2_lnot17_i1836 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv1_i_i1860_stall_local;
wire [63:0] local_bb2_conv1_i_i1860;

assign local_bb2_conv1_i_i1860[63:32] = 32'h0;
assign local_bb2_conv1_i_i1860[31:0] = local_bb2_or47_i1858;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot8_i1375_stall_local;
wire local_bb2_lnot8_i1375;

assign local_bb2_lnot8_i1375 = (local_bb2_and3_i1369 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_i1377_stall_local;
wire local_bb2_cmp11_i1377;

assign local_bb2_cmp11_i1377 = (local_bb2_and3_i1369 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u23_stall_local;
wire [31:0] local_bb2_var__u23;

assign local_bb2_var__u23 = (local_bb2_and3_i1369 | local_bb2_and6_i1373);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_not_i1383_stall_local;
wire local_bb2_lnot17_not_i1383;

assign local_bb2_lnot17_not_i1383 = (local_bb2_lnot17_i1379 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv1_i_i1403_stall_local;
wire [63:0] local_bb2_conv1_i_i1403;

assign local_bb2_conv1_i_i1403[63:32] = 32'h0;
assign local_bb2_conv1_i_i1403[31:0] = local_bb2_or47_i1401;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u24_stall_local;
wire [31:0] local_bb2_var__u24;

assign local_bb2_var__u24 = rnode_177to178_bb2_c0_ene5_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u25_stall_local;
wire [31:0] local_bb2_var__u25;

assign local_bb2_var__u25 = rnode_177to178_bb2_c0_ene6_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot8_i827_stall_local;
wire local_bb2_lnot8_i827;

assign local_bb2_lnot8_i827 = (local_bb2_and3_i821 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_i829_stall_local;
wire local_bb2_cmp11_i829;

assign local_bb2_cmp11_i829 = (local_bb2_and3_i821 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u26_stall_local;
wire [31:0] local_bb2_var__u26;

assign local_bb2_var__u26 = (local_bb2_and3_i821 | local_bb2_and6_i825);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_not_i835_stall_local;
wire local_bb2_lnot17_not_i835;

assign local_bb2_lnot17_not_i835 = (local_bb2_lnot17_i831 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv1_i_i855_stall_local;
wire [63:0] local_bb2_conv1_i_i855;

assign local_bb2_conv1_i_i855[63:32] = 32'h0;
assign local_bb2_conv1_i_i855[31:0] = local_bb2_or47_i853;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot8_i271_stall_local;
wire local_bb2_lnot8_i271;

assign local_bb2_lnot8_i271 = (local_bb2_and3_i265 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_i273_stall_local;
wire local_bb2_cmp11_i273;

assign local_bb2_cmp11_i273 = (local_bb2_and3_i265 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u27_stall_local;
wire [31:0] local_bb2_var__u27;

assign local_bb2_var__u27 = (local_bb2_and3_i265 | local_bb2_and6_i269);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_not_i279_stall_local;
wire local_bb2_lnot17_not_i279;

assign local_bb2_lnot17_not_i279 = (local_bb2_lnot17_i275 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv1_i_i299_stall_local;
wire [63:0] local_bb2_conv1_i_i299;

assign local_bb2_conv1_i_i299[63:32] = 32'h0;
assign local_bb2_conv1_i_i299[31:0] = local_bb2_or47_i297;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot8_i735_stall_local;
wire local_bb2_lnot8_i735;

assign local_bb2_lnot8_i735 = (local_bb2_and3_i729 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_i737_stall_local;
wire local_bb2_cmp11_i737;

assign local_bb2_cmp11_i737 = (local_bb2_and3_i729 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u28_stall_local;
wire [31:0] local_bb2_var__u28;

assign local_bb2_var__u28 = (local_bb2_and3_i729 | local_bb2_and6_i733);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_not_i743_stall_local;
wire local_bb2_lnot17_not_i743;

assign local_bb2_lnot17_not_i743 = (local_bb2_lnot17_i739 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv1_i_i763_stall_local;
wire [63:0] local_bb2_conv1_i_i763;

assign local_bb2_conv1_i_i763[63:32] = 32'h0;
assign local_bb2_conv1_i_i763[31:0] = local_bb2_or47_i761;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot8_i363_stall_local;
wire local_bb2_lnot8_i363;

assign local_bb2_lnot8_i363 = (local_bb2_and3_i357 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_i365_stall_local;
wire local_bb2_cmp11_i365;

assign local_bb2_cmp11_i365 = (local_bb2_and3_i357 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u29_stall_local;
wire [31:0] local_bb2_var__u29;

assign local_bb2_var__u29 = (local_bb2_and3_i357 | local_bb2_and6_i361);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot17_not_i371_stall_local;
wire local_bb2_lnot17_not_i371;

assign local_bb2_lnot17_not_i371 = (local_bb2_lnot17_i367 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv1_i_i391_stall_local;
wire [63:0] local_bb2_conv1_i_i391;

assign local_bb2_conv1_i_i391[63:32] = 32'h0;
assign local_bb2_conv1_i_i391[31:0] = local_bb2_or47_i389;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i_stall_local;
wire local_bb2_lnot_i;

assign local_bb2_lnot_i = (local_bb2_and_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i_stall_local;
wire local_bb2_cmp_i;

assign local_bb2_cmp_i = (local_bb2_and_i == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u30_stall_local;
wire [31:0] local_bb2_var__u30;

assign local_bb2_var__u30 = (local_bb2_and6_i | local_bb2_and_i);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i_stall_local;
wire [31:0] local_bb2_add_i;

assign local_bb2_add_i = (local_bb2_and3_i + local_bb2_and_i);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_not_i_stall_local;
wire local_bb2_lnot14_not_i;

assign local_bb2_lnot14_not_i = (local_bb2_lnot14_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv_i_i_stall_local;
wire [63:0] local_bb2_conv_i_i;

assign local_bb2_conv_i_i[63:32] = 32'h0;
assign local_bb2_conv_i_i[31:0] = local_bb2_or_i;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i1374_stall_local;
wire local_bb2_lnot_i1374;

assign local_bb2_lnot_i1374 = (local_bb2_and_i1367 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i1376_stall_local;
wire local_bb2_cmp_i1376;

assign local_bb2_cmp_i1376 = (local_bb2_and_i1367 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u31_stall_local;
wire [31:0] local_bb2_var__u31;

assign local_bb2_var__u31 = (local_bb2_and6_i1373 | local_bb2_and_i1367);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i1411_stall_local;
wire [31:0] local_bb2_add_i1411;

assign local_bb2_add_i1411 = (local_bb2_and3_i1369 + local_bb2_and_i1367);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_not_i1397_stall_local;
wire local_bb2_lnot14_not_i1397;

assign local_bb2_lnot14_not_i1397 = (local_bb2_lnot14_i1378 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv_i_i1402_stall_local;
wire [63:0] local_bb2_conv_i_i1402;

assign local_bb2_conv_i_i1402[63:32] = 32'h0;
assign local_bb2_conv_i_i1402[31:0] = local_bb2_or_i1400;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i826_stall_local;
wire local_bb2_lnot_i826;

assign local_bb2_lnot_i826 = (local_bb2_and_i819 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i828_stall_local;
wire local_bb2_cmp_i828;

assign local_bb2_cmp_i828 = (local_bb2_and_i819 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u32_stall_local;
wire [31:0] local_bb2_var__u32;

assign local_bb2_var__u32 = (local_bb2_and6_i825 | local_bb2_and_i819);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i863_stall_local;
wire [31:0] local_bb2_add_i863;

assign local_bb2_add_i863 = (local_bb2_and3_i821 + local_bb2_and_i819);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_not_i849_stall_local;
wire local_bb2_lnot14_not_i849;

assign local_bb2_lnot14_not_i849 = (local_bb2_lnot14_i830 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv_i_i854_stall_local;
wire [63:0] local_bb2_conv_i_i854;

assign local_bb2_conv_i_i854[63:32] = 32'h0;
assign local_bb2_conv_i_i854[31:0] = local_bb2_or_i852;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i362_stall_local;
wire local_bb2_lnot_i362;

assign local_bb2_lnot_i362 = (local_bb2_and_i355 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i364_stall_local;
wire local_bb2_cmp_i364;

assign local_bb2_cmp_i364 = (local_bb2_and_i355 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u33_stall_local;
wire [31:0] local_bb2_var__u33;

assign local_bb2_var__u33 = (local_bb2_and6_i361 | local_bb2_and_i355);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i399_stall_local;
wire [31:0] local_bb2_add_i399;

assign local_bb2_add_i399 = (local_bb2_and3_i357 + local_bb2_and_i355);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_not_i385_stall_local;
wire local_bb2_lnot14_not_i385;

assign local_bb2_lnot14_not_i385 = (local_bb2_lnot14_i366 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv_i_i390_stall_local;
wire [63:0] local_bb2_conv_i_i390;

assign local_bb2_conv_i_i390[63:32] = 32'h0;
assign local_bb2_conv_i_i390[31:0] = local_bb2_or_i388;

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge8_demorgan_i_stall_local;
wire local_bb2_brmerge8_demorgan_i;

assign local_bb2_brmerge8_demorgan_i = (local_bb2_cmp11_i & local_bb2_lnot17_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_not_i_stall_local;
wire local_bb2_cmp11_not_i;

assign local_bb2_cmp11_not_i = (local_bb2_cmp11_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u34_stall_local;
wire local_bb2_var__u34;

assign local_bb2_var__u34 = (local_bb2_var__u20 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge8_demorgan_i1288_stall_local;
wire local_bb2_brmerge8_demorgan_i1288;

assign local_bb2_brmerge8_demorgan_i1288 = (local_bb2_cmp11_i1285 & local_bb2_lnot17_i1287);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_not_i1292_stall_local;
wire local_bb2_cmp11_not_i1292;

assign local_bb2_cmp11_not_i1292 = (local_bb2_cmp11_i1285 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u35_stall_local;
wire local_bb2_var__u35;

assign local_bb2_var__u35 = (local_bb2_var__u21 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i1831_stall_local;
wire local_bb2_lnot_i1831;

assign local_bb2_lnot_i1831 = (local_bb2_and_i1824 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i1833_stall_local;
wire local_bb2_cmp_i1833;

assign local_bb2_cmp_i1833 = (local_bb2_and_i1824 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u36_stall_local;
wire [31:0] local_bb2_var__u36;

assign local_bb2_var__u36 = (local_bb2_and6_i1830 | local_bb2_and_i1824);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i1868_stall_local;
wire [31:0] local_bb2_add_i1868;

assign local_bb2_add_i1868 = (local_bb2_and3_i1826 + local_bb2_and_i1824);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_not_i1854_stall_local;
wire local_bb2_lnot14_not_i1854;

assign local_bb2_lnot14_not_i1854 = (local_bb2_lnot14_i1835 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv_i_i1859_stall_local;
wire [63:0] local_bb2_conv_i_i1859;

assign local_bb2_conv_i_i1859[63:32] = 32'h0;
assign local_bb2_conv_i_i1859[31:0] = local_bb2_or_i1857;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i1282_stall_local;
wire local_bb2_lnot_i1282;

assign local_bb2_lnot_i1282 = (local_bb2_and_i1275 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i1284_stall_local;
wire local_bb2_cmp_i1284;

assign local_bb2_cmp_i1284 = (local_bb2_and_i1275 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u37_stall_local;
wire [31:0] local_bb2_var__u37;

assign local_bb2_var__u37 = (local_bb2_and6_i1281 | local_bb2_and_i1275);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i1319_stall_local;
wire [31:0] local_bb2_add_i1319;

assign local_bb2_add_i1319 = (local_bb2_and3_i1277 + local_bb2_and_i1275);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_not_i1305_stall_local;
wire local_bb2_lnot14_not_i1305;

assign local_bb2_lnot14_not_i1305 = (local_bb2_lnot14_i1286 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv_i_i1310_stall_local;
wire [63:0] local_bb2_conv_i_i1310;

assign local_bb2_conv_i_i1310[63:32] = 32'h0;
assign local_bb2_conv_i_i1310[31:0] = local_bb2_or_i1308;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i734_stall_local;
wire local_bb2_lnot_i734;

assign local_bb2_lnot_i734 = (local_bb2_and_i727 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i736_stall_local;
wire local_bb2_cmp_i736;

assign local_bb2_cmp_i736 = (local_bb2_and_i727 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u38_stall_local;
wire [31:0] local_bb2_var__u38;

assign local_bb2_var__u38 = (local_bb2_and6_i733 | local_bb2_and_i727);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i771_stall_local;
wire [31:0] local_bb2_add_i771;

assign local_bb2_add_i771 = (local_bb2_and3_i729 + local_bb2_and_i727);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_not_i757_stall_local;
wire local_bb2_lnot14_not_i757;

assign local_bb2_lnot14_not_i757 = (local_bb2_lnot14_i738 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv_i_i762_stall_local;
wire [63:0] local_bb2_conv_i_i762;

assign local_bb2_conv_i_i762[63:32] = 32'h0;
assign local_bb2_conv_i_i762[31:0] = local_bb2_or_i760;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i270_stall_local;
wire local_bb2_lnot_i270;

assign local_bb2_lnot_i270 = (local_bb2_and_i263 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i272_stall_local;
wire local_bb2_cmp_i272;

assign local_bb2_cmp_i272 = (local_bb2_and_i263 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u39_stall_local;
wire [31:0] local_bb2_var__u39;

assign local_bb2_var__u39 = (local_bb2_and6_i269 | local_bb2_and_i263);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i307_stall_local;
wire [31:0] local_bb2_add_i307;

assign local_bb2_add_i307 = (local_bb2_and3_i265 + local_bb2_and_i263);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot14_not_i293_stall_local;
wire local_bb2_lnot14_not_i293;

assign local_bb2_lnot14_not_i293 = (local_bb2_lnot14_i274 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_conv_i_i298_stall_local;
wire [63:0] local_bb2_conv_i_i298;

assign local_bb2_conv_i_i298[63:32] = 32'h0;
assign local_bb2_conv_i_i298[31:0] = local_bb2_or_i296;

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge8_demorgan_i1837_stall_local;
wire local_bb2_brmerge8_demorgan_i1837;

assign local_bb2_brmerge8_demorgan_i1837 = (local_bb2_cmp11_i1834 & local_bb2_lnot17_i1836);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_not_i1841_stall_local;
wire local_bb2_cmp11_not_i1841;

assign local_bb2_cmp11_not_i1841 = (local_bb2_cmp11_i1834 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u40_stall_local;
wire local_bb2_var__u40;

assign local_bb2_var__u40 = (local_bb2_var__u22 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge8_demorgan_i1380_stall_local;
wire local_bb2_brmerge8_demorgan_i1380;

assign local_bb2_brmerge8_demorgan_i1380 = (local_bb2_cmp11_i1377 & local_bb2_lnot17_i1379);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_not_i1384_stall_local;
wire local_bb2_cmp11_not_i1384;

assign local_bb2_cmp11_not_i1384 = (local_bb2_cmp11_i1377 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u41_stall_local;
wire local_bb2_var__u41;

assign local_bb2_var__u41 = (local_bb2_var__u23 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_and2_i1460_stall_local;
wire [31:0] local_bb2_and2_i1460;

assign local_bb2_and2_i1460 = (local_bb2_var__u24 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and12_i1465_stall_local;
wire [31:0] local_bb2_and12_i1465;

assign local_bb2_and12_i1465 = (local_bb2_var__u24 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and2_i912_stall_local;
wire [31:0] local_bb2_and2_i912;

assign local_bb2_and2_i912 = (local_bb2_var__u25 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and12_i917_stall_local;
wire [31:0] local_bb2_and12_i917;

assign local_bb2_and12_i917 = (local_bb2_var__u25 & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge8_demorgan_i832_stall_local;
wire local_bb2_brmerge8_demorgan_i832;

assign local_bb2_brmerge8_demorgan_i832 = (local_bb2_cmp11_i829 & local_bb2_lnot17_i831);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_not_i836_stall_local;
wire local_bb2_cmp11_not_i836;

assign local_bb2_cmp11_not_i836 = (local_bb2_cmp11_i829 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u42_stall_local;
wire local_bb2_var__u42;

assign local_bb2_var__u42 = (local_bb2_var__u26 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge8_demorgan_i276_stall_local;
wire local_bb2_brmerge8_demorgan_i276;

assign local_bb2_brmerge8_demorgan_i276 = (local_bb2_cmp11_i273 & local_bb2_lnot17_i275);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_not_i280_stall_local;
wire local_bb2_cmp11_not_i280;

assign local_bb2_cmp11_not_i280 = (local_bb2_cmp11_i273 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u43_stall_local;
wire local_bb2_var__u43;

assign local_bb2_var__u43 = (local_bb2_var__u27 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge8_demorgan_i740_stall_local;
wire local_bb2_brmerge8_demorgan_i740;

assign local_bb2_brmerge8_demorgan_i740 = (local_bb2_cmp11_i737 & local_bb2_lnot17_i739);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_not_i744_stall_local;
wire local_bb2_cmp11_not_i744;

assign local_bb2_cmp11_not_i744 = (local_bb2_cmp11_i737 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u44_stall_local;
wire local_bb2_var__u44;

assign local_bb2_var__u44 = (local_bb2_var__u28 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge8_demorgan_i368_stall_local;
wire local_bb2_brmerge8_demorgan_i368;

assign local_bb2_brmerge8_demorgan_i368 = (local_bb2_cmp11_i365 & local_bb2_lnot17_i367);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp11_not_i372_stall_local;
wire local_bb2_cmp11_not_i372;

assign local_bb2_cmp11_not_i372 = (local_bb2_cmp11_i365 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u45_stall_local;
wire local_bb2_var__u45;

assign local_bb2_var__u45 = (local_bb2_var__u29 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i_stall_local;
wire local_bb2_reduction_0_i;

assign local_bb2_reduction_0_i = (local_bb2_lnot_i | local_bb2_lnot8_i);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u46_stall_local;
wire local_bb2_var__u46;

assign local_bb2_var__u46 = (local_bb2_cmp_i | local_bb2_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u47_stall_local;
wire local_bb2_var__u47;

assign local_bb2_var__u47 = (local_bb2_var__u30 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i_stall_local;
wire local_bb2__28_i;

assign local_bb2__28_i = (local_bb2_cmp_i & local_bb2_lnot14_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i1429_stall_local;
wire local_bb2_reduction_0_i1429;

assign local_bb2_reduction_0_i1429 = (local_bb2_lnot_i1374 | local_bb2_lnot8_i1375);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u48_stall_local;
wire local_bb2_var__u48;

assign local_bb2_var__u48 = (local_bb2_cmp_i1376 | local_bb2_cmp11_i1377);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u49_stall_local;
wire local_bb2_var__u49;

assign local_bb2_var__u49 = (local_bb2_var__u31 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i1398_stall_local;
wire local_bb2__28_i1398;

assign local_bb2__28_i1398 = (local_bb2_cmp_i1376 & local_bb2_lnot14_not_i1397);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i881_stall_local;
wire local_bb2_reduction_0_i881;

assign local_bb2_reduction_0_i881 = (local_bb2_lnot_i826 | local_bb2_lnot8_i827);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u50_stall_local;
wire local_bb2_var__u50;

assign local_bb2_var__u50 = (local_bb2_cmp_i828 | local_bb2_cmp11_i829);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u51_stall_local;
wire local_bb2_var__u51;

assign local_bb2_var__u51 = (local_bb2_var__u32 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i850_stall_local;
wire local_bb2__28_i850;

assign local_bb2__28_i850 = (local_bb2_cmp_i828 & local_bb2_lnot14_not_i849);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i417_stall_local;
wire local_bb2_reduction_0_i417;

assign local_bb2_reduction_0_i417 = (local_bb2_lnot_i362 | local_bb2_lnot8_i363);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u52_stall_local;
wire local_bb2_var__u52;

assign local_bb2_var__u52 = (local_bb2_cmp_i364 | local_bb2_cmp11_i365);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u53_stall_local;
wire local_bb2_var__u53;

assign local_bb2_var__u53 = (local_bb2_var__u33 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i386_stall_local;
wire local_bb2__28_i386;

assign local_bb2__28_i386 = (local_bb2_cmp_i364 & local_bb2_lnot14_not_i385);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge10_demorgan_i_stall_local;
wire local_bb2_brmerge10_demorgan_i;

assign local_bb2_brmerge10_demorgan_i = (local_bb2_brmerge8_demorgan_i & local_bb2_lnot_i);

// This section implements an unregistered operation.
// 
wire local_bb2__mux9_mux_i_stall_local;
wire local_bb2__mux9_mux_i;

assign local_bb2__mux9_mux_i = (local_bb2_brmerge8_demorgan_i ^ local_bb2_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge3_i_stall_local;
wire local_bb2_brmerge3_i;

assign local_bb2_brmerge3_i = (local_bb2_var__u34 | local_bb2_cmp11_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_i_stall_local;
wire local_bb2__mux_mux_i;

assign local_bb2__mux_mux_i = (local_bb2_var__u34 | local_bb2_cmp11_i);

// This section implements an unregistered operation.
// 
wire local_bb2__not_i_stall_local;
wire local_bb2__not_i;

assign local_bb2__not_i = (local_bb2_var__u34 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__mux9_mux_i1290_stall_local;
wire local_bb2__mux9_mux_i1290;

assign local_bb2__mux9_mux_i1290 = (local_bb2_brmerge8_demorgan_i1288 ^ local_bb2_cmp11_i1285);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge3_i1293_stall_local;
wire local_bb2_brmerge3_i1293;

assign local_bb2_brmerge3_i1293 = (local_bb2_var__u35 | local_bb2_cmp11_not_i1292);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_i1295_stall_local;
wire local_bb2__mux_mux_i1295;

assign local_bb2__mux_mux_i1295 = (local_bb2_var__u35 | local_bb2_cmp11_i1285);

// This section implements an unregistered operation.
// 
wire local_bb2__not_i1297_stall_local;
wire local_bb2__not_i1297;

assign local_bb2__not_i1297 = (local_bb2_var__u35 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i1886_stall_local;
wire local_bb2_reduction_0_i1886;

assign local_bb2_reduction_0_i1886 = (local_bb2_lnot_i1831 | local_bb2_lnot8_i1832);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u54_stall_local;
wire local_bb2_var__u54;

assign local_bb2_var__u54 = (local_bb2_cmp_i1833 | local_bb2_cmp11_i1834);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u55_stall_local;
wire local_bb2_var__u55;

assign local_bb2_var__u55 = (local_bb2_var__u36 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i1855_stall_local;
wire local_bb2__28_i1855;

assign local_bb2__28_i1855 = (local_bb2_cmp_i1833 & local_bb2_lnot14_not_i1854);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge10_demorgan_i1289_stall_local;
wire local_bb2_brmerge10_demorgan_i1289;

assign local_bb2_brmerge10_demorgan_i1289 = (local_bb2_brmerge8_demorgan_i1288 & local_bb2_lnot_i1282);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i1337_stall_local;
wire local_bb2_reduction_0_i1337;

assign local_bb2_reduction_0_i1337 = (local_bb2_lnot_i1282 | local_bb2_lnot8_i1283);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u56_stall_local;
wire local_bb2_var__u56;

assign local_bb2_var__u56 = (local_bb2_cmp_i1284 | local_bb2_cmp11_i1285);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u57_stall_local;
wire local_bb2_var__u57;

assign local_bb2_var__u57 = (local_bb2_var__u37 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i1306_stall_local;
wire local_bb2__28_i1306;

assign local_bb2__28_i1306 = (local_bb2_cmp_i1284 & local_bb2_lnot14_not_i1305);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i789_stall_local;
wire local_bb2_reduction_0_i789;

assign local_bb2_reduction_0_i789 = (local_bb2_lnot_i734 | local_bb2_lnot8_i735);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u58_stall_local;
wire local_bb2_var__u58;

assign local_bb2_var__u58 = (local_bb2_cmp_i736 | local_bb2_cmp11_i737);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u59_stall_local;
wire local_bb2_var__u59;

assign local_bb2_var__u59 = (local_bb2_var__u38 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i758_stall_local;
wire local_bb2__28_i758;

assign local_bb2__28_i758 = (local_bb2_cmp_i736 & local_bb2_lnot14_not_i757);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i325_stall_local;
wire local_bb2_reduction_0_i325;

assign local_bb2_reduction_0_i325 = (local_bb2_lnot_i270 | local_bb2_lnot8_i271);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u60_stall_local;
wire local_bb2_var__u60;

assign local_bb2_var__u60 = (local_bb2_cmp_i272 | local_bb2_cmp11_i273);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u61_stall_local;
wire local_bb2_var__u61;

assign local_bb2_var__u61 = (local_bb2_var__u39 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i294_stall_local;
wire local_bb2__28_i294;

assign local_bb2__28_i294 = (local_bb2_cmp_i272 & local_bb2_lnot14_not_i293);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge10_demorgan_i1838_stall_local;
wire local_bb2_brmerge10_demorgan_i1838;

assign local_bb2_brmerge10_demorgan_i1838 = (local_bb2_brmerge8_demorgan_i1837 & local_bb2_lnot_i1831);

// This section implements an unregistered operation.
// 
wire local_bb2__mux9_mux_i1839_stall_local;
wire local_bb2__mux9_mux_i1839;

assign local_bb2__mux9_mux_i1839 = (local_bb2_brmerge8_demorgan_i1837 ^ local_bb2_cmp11_i1834);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge3_i1842_stall_local;
wire local_bb2_brmerge3_i1842;

assign local_bb2_brmerge3_i1842 = (local_bb2_var__u40 | local_bb2_cmp11_not_i1841);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_i1844_stall_local;
wire local_bb2__mux_mux_i1844;

assign local_bb2__mux_mux_i1844 = (local_bb2_var__u40 | local_bb2_cmp11_i1834);

// This section implements an unregistered operation.
// 
wire local_bb2__not_i1846_stall_local;
wire local_bb2__not_i1846;

assign local_bb2__not_i1846 = (local_bb2_var__u40 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge10_demorgan_i1381_stall_local;
wire local_bb2_brmerge10_demorgan_i1381;

assign local_bb2_brmerge10_demorgan_i1381 = (local_bb2_brmerge8_demorgan_i1380 & local_bb2_lnot_i1374);

// This section implements an unregistered operation.
// 
wire local_bb2__mux9_mux_i1382_stall_local;
wire local_bb2__mux9_mux_i1382;

assign local_bb2__mux9_mux_i1382 = (local_bb2_brmerge8_demorgan_i1380 ^ local_bb2_cmp11_i1377);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge3_i1385_stall_local;
wire local_bb2_brmerge3_i1385;

assign local_bb2_brmerge3_i1385 = (local_bb2_var__u41 | local_bb2_cmp11_not_i1384);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_i1387_stall_local;
wire local_bb2__mux_mux_i1387;

assign local_bb2__mux_mux_i1387 = (local_bb2_var__u41 | local_bb2_cmp11_i1377);

// This section implements an unregistered operation.
// 
wire local_bb2__not_i1389_stall_local;
wire local_bb2__not_i1389;

assign local_bb2__not_i1389 = (local_bb2_var__u41 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i1461_stall_local;
wire [31:0] local_bb2_shr3_i1461;

assign local_bb2_shr3_i1461 = (local_bb2_and2_i1460 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i913_stall_local;
wire [31:0] local_bb2_shr3_i913;

assign local_bb2_shr3_i913 = (local_bb2_and2_i912 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge10_demorgan_i833_stall_local;
wire local_bb2_brmerge10_demorgan_i833;

assign local_bb2_brmerge10_demorgan_i833 = (local_bb2_brmerge8_demorgan_i832 & local_bb2_lnot_i826);

// This section implements an unregistered operation.
// 
wire local_bb2__mux9_mux_i834_stall_local;
wire local_bb2__mux9_mux_i834;

assign local_bb2__mux9_mux_i834 = (local_bb2_brmerge8_demorgan_i832 ^ local_bb2_cmp11_i829);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge3_i837_stall_local;
wire local_bb2_brmerge3_i837;

assign local_bb2_brmerge3_i837 = (local_bb2_var__u42 | local_bb2_cmp11_not_i836);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_i839_stall_local;
wire local_bb2__mux_mux_i839;

assign local_bb2__mux_mux_i839 = (local_bb2_var__u42 | local_bb2_cmp11_i829);

// This section implements an unregistered operation.
// 
wire local_bb2__not_i841_stall_local;
wire local_bb2__not_i841;

assign local_bb2__not_i841 = (local_bb2_var__u42 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge10_demorgan_i277_stall_local;
wire local_bb2_brmerge10_demorgan_i277;

assign local_bb2_brmerge10_demorgan_i277 = (local_bb2_brmerge8_demorgan_i276 & local_bb2_lnot_i270);

// This section implements an unregistered operation.
// 
wire local_bb2__mux9_mux_i278_stall_local;
wire local_bb2__mux9_mux_i278;

assign local_bb2__mux9_mux_i278 = (local_bb2_brmerge8_demorgan_i276 ^ local_bb2_cmp11_i273);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge3_i281_stall_local;
wire local_bb2_brmerge3_i281;

assign local_bb2_brmerge3_i281 = (local_bb2_var__u43 | local_bb2_cmp11_not_i280);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_i283_stall_local;
wire local_bb2__mux_mux_i283;

assign local_bb2__mux_mux_i283 = (local_bb2_var__u43 | local_bb2_cmp11_i273);

// This section implements an unregistered operation.
// 
wire local_bb2__not_i285_stall_local;
wire local_bb2__not_i285;

assign local_bb2__not_i285 = (local_bb2_var__u43 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge10_demorgan_i741_stall_local;
wire local_bb2_brmerge10_demorgan_i741;

assign local_bb2_brmerge10_demorgan_i741 = (local_bb2_brmerge8_demorgan_i740 & local_bb2_lnot_i734);

// This section implements an unregistered operation.
// 
wire local_bb2__mux9_mux_i742_stall_local;
wire local_bb2__mux9_mux_i742;

assign local_bb2__mux9_mux_i742 = (local_bb2_brmerge8_demorgan_i740 ^ local_bb2_cmp11_i737);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge3_i745_stall_local;
wire local_bb2_brmerge3_i745;

assign local_bb2_brmerge3_i745 = (local_bb2_var__u44 | local_bb2_cmp11_not_i744);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_i747_stall_local;
wire local_bb2__mux_mux_i747;

assign local_bb2__mux_mux_i747 = (local_bb2_var__u44 | local_bb2_cmp11_i737);

// This section implements an unregistered operation.
// 
wire local_bb2__not_i749_stall_local;
wire local_bb2__not_i749;

assign local_bb2__not_i749 = (local_bb2_var__u44 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge10_demorgan_i369_stall_local;
wire local_bb2_brmerge10_demorgan_i369;

assign local_bb2_brmerge10_demorgan_i369 = (local_bb2_brmerge8_demorgan_i368 & local_bb2_lnot_i362);

// This section implements an unregistered operation.
// 
wire local_bb2__mux9_mux_i370_stall_local;
wire local_bb2__mux9_mux_i370;

assign local_bb2__mux9_mux_i370 = (local_bb2_brmerge8_demorgan_i368 ^ local_bb2_cmp11_i365);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge3_i373_stall_local;
wire local_bb2_brmerge3_i373;

assign local_bb2_brmerge3_i373 = (local_bb2_var__u45 | local_bb2_cmp11_not_i372);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_i375_stall_local;
wire local_bb2__mux_mux_i375;

assign local_bb2__mux_mux_i375 = (local_bb2_var__u45 | local_bb2_cmp11_i365);

// This section implements an unregistered operation.
// 
wire local_bb2__not_i377_stall_local;
wire local_bb2__not_i377;

assign local_bb2__not_i377 = (local_bb2_var__u45 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__26_demorgan_i_stall_local;
wire local_bb2__26_demorgan_i;

assign local_bb2__26_demorgan_i = (local_bb2_cmp_i | local_bb2_brmerge10_demorgan_i);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge5_i_stall_local;
wire local_bb2_brmerge5_i;

assign local_bb2_brmerge5_i = (local_bb2_brmerge3_i | local_bb2_lnot17_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i_stall_local;
wire local_bb2_reduction_3_i;

assign local_bb2_reduction_3_i = (local_bb2_cmp11_i & local_bb2__not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge5_i1294_stall_local;
wire local_bb2_brmerge5_i1294;

assign local_bb2_brmerge5_i1294 = (local_bb2_brmerge3_i1293 | local_bb2_lnot17_not_i1291);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i1298_stall_local;
wire local_bb2_reduction_3_i1298;

assign local_bb2_reduction_3_i1298 = (local_bb2_cmp11_i1285 & local_bb2__not_i1297);

// This section implements an unregistered operation.
// 
wire local_bb2__26_demorgan_i1303_stall_local;
wire local_bb2__26_demorgan_i1303;

assign local_bb2__26_demorgan_i1303 = (local_bb2_cmp_i1284 | local_bb2_brmerge10_demorgan_i1289);

// This section implements an unregistered operation.
// 
wire local_bb2__26_demorgan_i1852_stall_local;
wire local_bb2__26_demorgan_i1852;

assign local_bb2__26_demorgan_i1852 = (local_bb2_cmp_i1833 | local_bb2_brmerge10_demorgan_i1838);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge5_i1843_stall_local;
wire local_bb2_brmerge5_i1843;

assign local_bb2_brmerge5_i1843 = (local_bb2_brmerge3_i1842 | local_bb2_lnot17_not_i1840);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i1847_stall_local;
wire local_bb2_reduction_3_i1847;

assign local_bb2_reduction_3_i1847 = (local_bb2_cmp11_i1834 & local_bb2__not_i1846);

// This section implements an unregistered operation.
// 
wire local_bb2__26_demorgan_i1395_stall_local;
wire local_bb2__26_demorgan_i1395;

assign local_bb2__26_demorgan_i1395 = (local_bb2_cmp_i1376 | local_bb2_brmerge10_demorgan_i1381);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge5_i1386_stall_local;
wire local_bb2_brmerge5_i1386;

assign local_bb2_brmerge5_i1386 = (local_bb2_brmerge3_i1385 | local_bb2_lnot17_not_i1383);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i1390_stall_local;
wire local_bb2_reduction_3_i1390;

assign local_bb2_reduction_3_i1390 = (local_bb2_cmp11_i1377 & local_bb2__not_i1389);

// This section implements an unregistered operation.
// 
wire local_bb2__26_demorgan_i847_stall_local;
wire local_bb2__26_demorgan_i847;

assign local_bb2__26_demorgan_i847 = (local_bb2_cmp_i828 | local_bb2_brmerge10_demorgan_i833);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge5_i838_stall_local;
wire local_bb2_brmerge5_i838;

assign local_bb2_brmerge5_i838 = (local_bb2_brmerge3_i837 | local_bb2_lnot17_not_i835);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i842_stall_local;
wire local_bb2_reduction_3_i842;

assign local_bb2_reduction_3_i842 = (local_bb2_cmp11_i829 & local_bb2__not_i841);

// This section implements an unregistered operation.
// 
wire local_bb2__26_demorgan_i291_stall_local;
wire local_bb2__26_demorgan_i291;

assign local_bb2__26_demorgan_i291 = (local_bb2_cmp_i272 | local_bb2_brmerge10_demorgan_i277);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge5_i282_stall_local;
wire local_bb2_brmerge5_i282;

assign local_bb2_brmerge5_i282 = (local_bb2_brmerge3_i281 | local_bb2_lnot17_not_i279);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i286_stall_local;
wire local_bb2_reduction_3_i286;

assign local_bb2_reduction_3_i286 = (local_bb2_cmp11_i273 & local_bb2__not_i285);

// This section implements an unregistered operation.
// 
wire local_bb2__26_demorgan_i755_stall_local;
wire local_bb2__26_demorgan_i755;

assign local_bb2__26_demorgan_i755 = (local_bb2_cmp_i736 | local_bb2_brmerge10_demorgan_i741);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge5_i746_stall_local;
wire local_bb2_brmerge5_i746;

assign local_bb2_brmerge5_i746 = (local_bb2_brmerge3_i745 | local_bb2_lnot17_not_i743);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i750_stall_local;
wire local_bb2_reduction_3_i750;

assign local_bb2_reduction_3_i750 = (local_bb2_cmp11_i737 & local_bb2__not_i749);

// This section implements an unregistered operation.
// 
wire local_bb2__26_demorgan_i383_stall_local;
wire local_bb2__26_demorgan_i383;

assign local_bb2__26_demorgan_i383 = (local_bb2_cmp_i364 | local_bb2_brmerge10_demorgan_i369);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge5_i374_stall_local;
wire local_bb2_brmerge5_i374;

assign local_bb2_brmerge5_i374 = (local_bb2_brmerge3_i373 | local_bb2_lnot17_not_i371);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i378_stall_local;
wire local_bb2_reduction_3_i378;

assign local_bb2_reduction_3_i378 = (local_bb2_cmp11_i365 & local_bb2__not_i377);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_mux_i_stall_local;
wire local_bb2__mux_mux_mux_i;

assign local_bb2__mux_mux_mux_i = (local_bb2_brmerge5_i & local_bb2__mux_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i_stall_local;
wire local_bb2_reduction_5_i;

assign local_bb2_reduction_5_i = (local_bb2_lnot14_i & local_bb2_reduction_3_i);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_mux_i1296_stall_local;
wire local_bb2__mux_mux_mux_i1296;

assign local_bb2__mux_mux_mux_i1296 = (local_bb2_brmerge5_i1294 & local_bb2__mux_mux_i1295);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i1299_stall_local;
wire local_bb2_reduction_5_i1299;

assign local_bb2_reduction_5_i1299 = (local_bb2_lnot14_i1286 & local_bb2_reduction_3_i1298);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_mux_i1845_stall_local;
wire local_bb2__mux_mux_mux_i1845;

assign local_bb2__mux_mux_mux_i1845 = (local_bb2_brmerge5_i1843 & local_bb2__mux_mux_i1844);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i1848_stall_local;
wire local_bb2_reduction_5_i1848;

assign local_bb2_reduction_5_i1848 = (local_bb2_lnot14_i1835 & local_bb2_reduction_3_i1847);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_mux_i1388_stall_local;
wire local_bb2__mux_mux_mux_i1388;

assign local_bb2__mux_mux_mux_i1388 = (local_bb2_brmerge5_i1386 & local_bb2__mux_mux_i1387);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i1391_stall_local;
wire local_bb2_reduction_5_i1391;

assign local_bb2_reduction_5_i1391 = (local_bb2_lnot14_i1378 & local_bb2_reduction_3_i1390);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_mux_i840_stall_local;
wire local_bb2__mux_mux_mux_i840;

assign local_bb2__mux_mux_mux_i840 = (local_bb2_brmerge5_i838 & local_bb2__mux_mux_i839);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i843_stall_local;
wire local_bb2_reduction_5_i843;

assign local_bb2_reduction_5_i843 = (local_bb2_lnot14_i830 & local_bb2_reduction_3_i842);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_mux_i284_stall_local;
wire local_bb2__mux_mux_mux_i284;

assign local_bb2__mux_mux_mux_i284 = (local_bb2_brmerge5_i282 & local_bb2__mux_mux_i283);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i287_stall_local;
wire local_bb2_reduction_5_i287;

assign local_bb2_reduction_5_i287 = (local_bb2_lnot14_i274 & local_bb2_reduction_3_i286);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_mux_i748_stall_local;
wire local_bb2__mux_mux_mux_i748;

assign local_bb2__mux_mux_mux_i748 = (local_bb2_brmerge5_i746 & local_bb2__mux_mux_i747);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i751_stall_local;
wire local_bb2_reduction_5_i751;

assign local_bb2_reduction_5_i751 = (local_bb2_lnot14_i738 & local_bb2_reduction_3_i750);

// This section implements an unregistered operation.
// 
wire local_bb2__mux_mux_mux_i376_stall_local;
wire local_bb2__mux_mux_mux_i376;

assign local_bb2__mux_mux_mux_i376 = (local_bb2_brmerge5_i374 & local_bb2__mux_mux_i375);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i379_stall_local;
wire local_bb2_reduction_5_i379;

assign local_bb2_reduction_5_i379 = (local_bb2_lnot14_i366 & local_bb2_reduction_3_i378);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i_stall_local;
wire local_bb2_reduction_6_i;

assign local_bb2_reduction_6_i = (local_bb2_var__u47 & local_bb2_reduction_5_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i1300_stall_local;
wire local_bb2_reduction_6_i1300;

assign local_bb2_reduction_6_i1300 = (local_bb2_var__u57 & local_bb2_reduction_5_i1299);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i1849_stall_local;
wire local_bb2_reduction_6_i1849;

assign local_bb2_reduction_6_i1849 = (local_bb2_var__u55 & local_bb2_reduction_5_i1848);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i1392_stall_local;
wire local_bb2_reduction_6_i1392;

assign local_bb2_reduction_6_i1392 = (local_bb2_var__u49 & local_bb2_reduction_5_i1391);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i844_stall_local;
wire local_bb2_reduction_6_i844;

assign local_bb2_reduction_6_i844 = (local_bb2_var__u51 & local_bb2_reduction_5_i843);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i288_stall_local;
wire local_bb2_reduction_6_i288;

assign local_bb2_reduction_6_i288 = (local_bb2_var__u61 & local_bb2_reduction_5_i287);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i752_stall_local;
wire local_bb2_reduction_6_i752;

assign local_bb2_reduction_6_i752 = (local_bb2_var__u59 & local_bb2_reduction_5_i751);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i380_stall_local;
wire local_bb2_reduction_6_i380;

assign local_bb2_reduction_6_i380 = (local_bb2_var__u53 & local_bb2_reduction_5_i379);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i_stall_local;
wire local_bb2__24_i;

assign local_bb2__24_i = (local_bb2_cmp_i ? local_bb2_reduction_6_i : local_bb2_brmerge10_demorgan_i);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i1301_stall_local;
wire local_bb2__24_i1301;

assign local_bb2__24_i1301 = (local_bb2_cmp_i1284 ? local_bb2_reduction_6_i1300 : local_bb2_brmerge10_demorgan_i1289);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i1850_stall_local;
wire local_bb2__24_i1850;

assign local_bb2__24_i1850 = (local_bb2_cmp_i1833 ? local_bb2_reduction_6_i1849 : local_bb2_brmerge10_demorgan_i1838);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i1393_stall_local;
wire local_bb2__24_i1393;

assign local_bb2__24_i1393 = (local_bb2_cmp_i1376 ? local_bb2_reduction_6_i1392 : local_bb2_brmerge10_demorgan_i1381);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i845_stall_local;
wire local_bb2__24_i845;

assign local_bb2__24_i845 = (local_bb2_cmp_i828 ? local_bb2_reduction_6_i844 : local_bb2_brmerge10_demorgan_i833);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i289_stall_local;
wire local_bb2__24_i289;

assign local_bb2__24_i289 = (local_bb2_cmp_i272 ? local_bb2_reduction_6_i288 : local_bb2_brmerge10_demorgan_i277);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i753_stall_local;
wire local_bb2__24_i753;

assign local_bb2__24_i753 = (local_bb2_cmp_i736 ? local_bb2_reduction_6_i752 : local_bb2_brmerge10_demorgan_i741);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i381_stall_local;
wire local_bb2__24_i381;

assign local_bb2__24_i381 = (local_bb2_cmp_i364 ? local_bb2_reduction_6_i380 : local_bb2_brmerge10_demorgan_i369);

// This section implements an unregistered operation.
// 
wire local_bb2__25_i_stall_local;
wire local_bb2__25_i;

assign local_bb2__25_i = (local_bb2__24_i ? local_bb2_lnot14_i : local_bb2__mux_mux_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb2__25_i1302_stall_local;
wire local_bb2__25_i1302;

assign local_bb2__25_i1302 = (local_bb2__24_i1301 ? local_bb2_lnot14_i1286 : local_bb2__mux_mux_mux_i1296);

// This section implements an unregistered operation.
// 
wire local_bb2__25_i1851_stall_local;
wire local_bb2__25_i1851;

assign local_bb2__25_i1851 = (local_bb2__24_i1850 ? local_bb2_lnot14_i1835 : local_bb2__mux_mux_mux_i1845);

// This section implements an unregistered operation.
// 
wire local_bb2__25_i1394_stall_local;
wire local_bb2__25_i1394;

assign local_bb2__25_i1394 = (local_bb2__24_i1393 ? local_bb2_lnot14_i1378 : local_bb2__mux_mux_mux_i1388);

// This section implements an unregistered operation.
// 
wire local_bb2__25_i846_stall_local;
wire local_bb2__25_i846;

assign local_bb2__25_i846 = (local_bb2__24_i845 ? local_bb2_lnot14_i830 : local_bb2__mux_mux_mux_i840);

// This section implements an unregistered operation.
// 
wire local_bb2__25_i290_stall_local;
wire local_bb2__25_i290;

assign local_bb2__25_i290 = (local_bb2__24_i289 ? local_bb2_lnot14_i274 : local_bb2__mux_mux_mux_i284);

// This section implements an unregistered operation.
// 
wire local_bb2__25_i754_stall_local;
wire local_bb2__25_i754;

assign local_bb2__25_i754 = (local_bb2__24_i753 ? local_bb2_lnot14_i738 : local_bb2__mux_mux_mux_i748);

// This section implements an unregistered operation.
// 
wire local_bb2__25_i382_stall_local;
wire local_bb2__25_i382;

assign local_bb2__25_i382 = (local_bb2__24_i381 ? local_bb2_lnot14_i366 : local_bb2__mux_mux_mux_i376);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i_stall_local;
wire local_bb2__27_i;

assign local_bb2__27_i = (local_bb2__26_demorgan_i ? local_bb2__25_i : local_bb2__mux9_mux_i);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i1304_stall_local;
wire local_bb2__27_i1304;

assign local_bb2__27_i1304 = (local_bb2__26_demorgan_i1303 ? local_bb2__25_i1302 : local_bb2__mux9_mux_i1290);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i1853_stall_local;
wire local_bb2__27_i1853;

assign local_bb2__27_i1853 = (local_bb2__26_demorgan_i1852 ? local_bb2__25_i1851 : local_bb2__mux9_mux_i1839);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i1396_stall_local;
wire local_bb2__27_i1396;

assign local_bb2__27_i1396 = (local_bb2__26_demorgan_i1395 ? local_bb2__25_i1394 : local_bb2__mux9_mux_i1382);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i848_stall_local;
wire local_bb2__27_i848;

assign local_bb2__27_i848 = (local_bb2__26_demorgan_i847 ? local_bb2__25_i846 : local_bb2__mux9_mux_i834);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i292_stall_local;
wire local_bb2__27_i292;

assign local_bb2__27_i292 = (local_bb2__26_demorgan_i291 ? local_bb2__25_i290 : local_bb2__mux9_mux_i278);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i756_stall_local;
wire local_bb2__27_i756;

assign local_bb2__27_i756 = (local_bb2__26_demorgan_i755 ? local_bb2__25_i754 : local_bb2__mux9_mux_i742);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i384_stall_local;
wire local_bb2__27_i384;

assign local_bb2__27_i384 = (local_bb2__26_demorgan_i383 ? local_bb2__25_i382 : local_bb2__mux9_mux_i370);

// This section implements an unregistered operation.
// 
wire local_bb2__29_i_stall_local;
wire local_bb2__29_i;

assign local_bb2__29_i = (local_bb2__28_i | local_bb2__27_i);

// This section implements an unregistered operation.
// 
wire local_bb2__29_i1307_stall_local;
wire local_bb2__29_i1307;

assign local_bb2__29_i1307 = (local_bb2__28_i1306 | local_bb2__27_i1304);

// This section implements an unregistered operation.
// 
wire local_bb2__29_i1856_stall_local;
wire local_bb2__29_i1856;

assign local_bb2__29_i1856 = (local_bb2__28_i1855 | local_bb2__27_i1853);

// This section implements an unregistered operation.
// 
wire local_bb2__29_i1399_stall_local;
wire local_bb2__29_i1399;

assign local_bb2__29_i1399 = (local_bb2__28_i1398 | local_bb2__27_i1396);

// This section implements an unregistered operation.
// 
wire local_bb2__29_i851_stall_local;
wire local_bb2__29_i851;

assign local_bb2__29_i851 = (local_bb2__28_i850 | local_bb2__27_i848);

// This section implements an unregistered operation.
// 
wire local_bb2__29_i295_stall_local;
wire local_bb2__29_i295;

assign local_bb2__29_i295 = (local_bb2__28_i294 | local_bb2__27_i292);

// This section implements an unregistered operation.
// 
wire local_bb2__29_i759_stall_local;
wire local_bb2__29_i759;

assign local_bb2__29_i759 = (local_bb2__28_i758 | local_bb2__27_i756);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i_valid_out;
wire local_bb2_xor_i_stall_in;
 reg local_bb2_xor_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_xor_i1278_valid_out;
wire local_bb2_xor_i1278_stall_in;
 reg local_bb2_xor_i1278_consumed_0_NO_SHIFT_REG;
wire local_bb2_xor_i1827_valid_out;
wire local_bb2_xor_i1827_stall_in;
 reg local_bb2_xor_i1827_consumed_0_NO_SHIFT_REG;
wire local_bb2_xor_i1370_valid_out;
wire local_bb2_xor_i1370_stall_in;
 reg local_bb2_xor_i1370_consumed_0_NO_SHIFT_REG;
wire local_bb2_xor_i822_valid_out;
wire local_bb2_xor_i822_stall_in;
 reg local_bb2_xor_i822_consumed_0_NO_SHIFT_REG;
wire local_bb2_xor_i266_valid_out;
wire local_bb2_xor_i266_stall_in;
 reg local_bb2_xor_i266_consumed_0_NO_SHIFT_REG;
wire local_bb2_xor_i730_valid_out;
wire local_bb2_xor_i730_stall_in;
 reg local_bb2_xor_i730_consumed_0_NO_SHIFT_REG;
wire local_bb2_xor_i358_valid_out;
wire local_bb2_xor_i358_stall_in;
 reg local_bb2_xor_i358_consumed_0_NO_SHIFT_REG;
wire local_bb2_add_i_valid_out;
wire local_bb2_add_i_stall_in;
 reg local_bb2_add_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv1_i_i_valid_out;
wire local_bb2_conv1_i_i_stall_in;
 reg local_bb2_conv1_i_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_add_i1319_valid_out;
wire local_bb2_add_i1319_stall_in;
 reg local_bb2_add_i1319_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv1_i_i1311_valid_out;
wire local_bb2_conv1_i_i1311_stall_in;
 reg local_bb2_conv1_i_i1311_consumed_0_NO_SHIFT_REG;
wire local_bb2_add_i1868_valid_out;
wire local_bb2_add_i1868_stall_in;
 reg local_bb2_add_i1868_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv1_i_i1860_valid_out;
wire local_bb2_conv1_i_i1860_stall_in;
 reg local_bb2_conv1_i_i1860_consumed_0_NO_SHIFT_REG;
wire local_bb2_add_i1411_valid_out;
wire local_bb2_add_i1411_stall_in;
 reg local_bb2_add_i1411_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv1_i_i1403_valid_out;
wire local_bb2_conv1_i_i1403_stall_in;
 reg local_bb2_conv1_i_i1403_consumed_0_NO_SHIFT_REG;
wire local_bb2_add_i863_valid_out;
wire local_bb2_add_i863_stall_in;
 reg local_bb2_add_i863_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv1_i_i855_valid_out;
wire local_bb2_conv1_i_i855_stall_in;
 reg local_bb2_conv1_i_i855_consumed_0_NO_SHIFT_REG;
wire local_bb2_add_i307_valid_out;
wire local_bb2_add_i307_stall_in;
 reg local_bb2_add_i307_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv1_i_i299_valid_out;
wire local_bb2_conv1_i_i299_stall_in;
 reg local_bb2_conv1_i_i299_consumed_0_NO_SHIFT_REG;
wire local_bb2_add_i771_valid_out;
wire local_bb2_add_i771_stall_in;
 reg local_bb2_add_i771_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv1_i_i763_valid_out;
wire local_bb2_conv1_i_i763_stall_in;
 reg local_bb2_conv1_i_i763_consumed_0_NO_SHIFT_REG;
wire local_bb2_add_i399_valid_out;
wire local_bb2_add_i399_stall_in;
 reg local_bb2_add_i399_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv1_i_i391_valid_out;
wire local_bb2_conv1_i_i391_stall_in;
 reg local_bb2_conv1_i_i391_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv_i_i_valid_out;
wire local_bb2_conv_i_i_stall_in;
 reg local_bb2_conv_i_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv_i_i1402_valid_out;
wire local_bb2_conv_i_i1402_stall_in;
 reg local_bb2_conv_i_i1402_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv_i_i854_valid_out;
wire local_bb2_conv_i_i854_stall_in;
 reg local_bb2_conv_i_i854_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv_i_i390_valid_out;
wire local_bb2_conv_i_i390_stall_in;
 reg local_bb2_conv_i_i390_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i_valid_out;
wire local_bb2_reduction_0_i_stall_in;
 reg local_bb2_reduction_0_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u46_valid_out;
wire local_bb2_var__u46_stall_in;
 reg local_bb2_var__u46_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i1337_valid_out;
wire local_bb2_reduction_0_i1337_stall_in;
 reg local_bb2_reduction_0_i1337_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u56_valid_out;
wire local_bb2_var__u56_stall_in;
 reg local_bb2_var__u56_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv_i_i1859_valid_out;
wire local_bb2_conv_i_i1859_stall_in;
 reg local_bb2_conv_i_i1859_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv_i_i1310_valid_out;
wire local_bb2_conv_i_i1310_stall_in;
 reg local_bb2_conv_i_i1310_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv_i_i762_valid_out;
wire local_bb2_conv_i_i762_stall_in;
 reg local_bb2_conv_i_i762_consumed_0_NO_SHIFT_REG;
wire local_bb2_conv_i_i298_valid_out;
wire local_bb2_conv_i_i298_stall_in;
 reg local_bb2_conv_i_i298_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i1886_valid_out;
wire local_bb2_reduction_0_i1886_stall_in;
 reg local_bb2_reduction_0_i1886_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u54_valid_out;
wire local_bb2_var__u54_stall_in;
 reg local_bb2_var__u54_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i1429_valid_out;
wire local_bb2_reduction_0_i1429_stall_in;
 reg local_bb2_reduction_0_i1429_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u48_valid_out;
wire local_bb2_var__u48_stall_in;
 reg local_bb2_var__u48_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i881_valid_out;
wire local_bb2_reduction_0_i881_stall_in;
 reg local_bb2_reduction_0_i881_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u50_valid_out;
wire local_bb2_var__u50_stall_in;
 reg local_bb2_var__u50_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i325_valid_out;
wire local_bb2_reduction_0_i325_stall_in;
 reg local_bb2_reduction_0_i325_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u60_valid_out;
wire local_bb2_var__u60_stall_in;
 reg local_bb2_var__u60_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i789_valid_out;
wire local_bb2_reduction_0_i789_stall_in;
 reg local_bb2_reduction_0_i789_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u58_valid_out;
wire local_bb2_var__u58_stall_in;
 reg local_bb2_var__u58_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i417_valid_out;
wire local_bb2_reduction_0_i417_stall_in;
 reg local_bb2_reduction_0_i417_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u52_valid_out;
wire local_bb2_var__u52_stall_in;
 reg local_bb2_var__u52_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i_valid_out;
wire local_bb2__29_i_stall_in;
 reg local_bb2__29_i_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i1399_valid_out;
wire local_bb2__29_i1399_stall_in;
 reg local_bb2__29_i1399_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i851_valid_out;
wire local_bb2__29_i851_stall_in;
 reg local_bb2__29_i851_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i387_valid_out;
wire local_bb2__29_i387_stall_in;
 reg local_bb2__29_i387_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i1307_valid_out;
wire local_bb2__29_i1307_stall_in;
 reg local_bb2__29_i1307_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i1856_valid_out;
wire local_bb2__29_i1856_stall_in;
 reg local_bb2__29_i1856_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i759_valid_out;
wire local_bb2__29_i759_stall_in;
 reg local_bb2__29_i759_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i295_valid_out;
wire local_bb2__29_i295_stall_in;
 reg local_bb2__29_i295_consumed_0_NO_SHIFT_REG;
wire local_bb2__29_i387_inputs_ready;
wire local_bb2__29_i387_stall_local;
wire local_bb2__29_i387;

assign local_bb2__29_i387_inputs_ready = (local_bb2_c0_enter_c0_eni8_valid_out_0_NO_SHIFT_REG & local_bb2_c0_enter_c0_eni8_valid_out_1_NO_SHIFT_REG & local_bb2_c0_enter_c0_eni8_valid_out_3_NO_SHIFT_REG & local_bb2_c0_enter_c0_eni8_valid_out_6_NO_SHIFT_REG & local_bb2_c0_enter_c0_eni8_valid_out_7_NO_SHIFT_REG & local_bb2_c0_enter_c0_eni8_valid_out_2_NO_SHIFT_REG);
assign local_bb2__29_i387 = (local_bb2__28_i386 | local_bb2__27_i384);
assign local_bb2_xor_i_valid_out = 1'b1;
assign local_bb2_xor_i1278_valid_out = 1'b1;
assign local_bb2_xor_i1827_valid_out = 1'b1;
assign local_bb2_xor_i1370_valid_out = 1'b1;
assign local_bb2_xor_i822_valid_out = 1'b1;
assign local_bb2_xor_i266_valid_out = 1'b1;
assign local_bb2_xor_i730_valid_out = 1'b1;
assign local_bb2_xor_i358_valid_out = 1'b1;
assign local_bb2_add_i_valid_out = 1'b1;
assign local_bb2_conv1_i_i_valid_out = 1'b1;
assign local_bb2_add_i1319_valid_out = 1'b1;
assign local_bb2_conv1_i_i1311_valid_out = 1'b1;
assign local_bb2_add_i1868_valid_out = 1'b1;
assign local_bb2_conv1_i_i1860_valid_out = 1'b1;
assign local_bb2_add_i1411_valid_out = 1'b1;
assign local_bb2_conv1_i_i1403_valid_out = 1'b1;
assign local_bb2_add_i863_valid_out = 1'b1;
assign local_bb2_conv1_i_i855_valid_out = 1'b1;
assign local_bb2_add_i307_valid_out = 1'b1;
assign local_bb2_conv1_i_i299_valid_out = 1'b1;
assign local_bb2_add_i771_valid_out = 1'b1;
assign local_bb2_conv1_i_i763_valid_out = 1'b1;
assign local_bb2_add_i399_valid_out = 1'b1;
assign local_bb2_conv1_i_i391_valid_out = 1'b1;
assign local_bb2_conv_i_i_valid_out = 1'b1;
assign local_bb2_conv_i_i1402_valid_out = 1'b1;
assign local_bb2_conv_i_i854_valid_out = 1'b1;
assign local_bb2_conv_i_i390_valid_out = 1'b1;
assign local_bb2_reduction_0_i_valid_out = 1'b1;
assign local_bb2_var__u46_valid_out = 1'b1;
assign local_bb2_reduction_0_i1337_valid_out = 1'b1;
assign local_bb2_var__u56_valid_out = 1'b1;
assign local_bb2_conv_i_i1859_valid_out = 1'b1;
assign local_bb2_conv_i_i1310_valid_out = 1'b1;
assign local_bb2_conv_i_i762_valid_out = 1'b1;
assign local_bb2_conv_i_i298_valid_out = 1'b1;
assign local_bb2_reduction_0_i1886_valid_out = 1'b1;
assign local_bb2_var__u54_valid_out = 1'b1;
assign local_bb2_reduction_0_i1429_valid_out = 1'b1;
assign local_bb2_var__u48_valid_out = 1'b1;
assign local_bb2_reduction_0_i881_valid_out = 1'b1;
assign local_bb2_var__u50_valid_out = 1'b1;
assign local_bb2_reduction_0_i325_valid_out = 1'b1;
assign local_bb2_var__u60_valid_out = 1'b1;
assign local_bb2_reduction_0_i789_valid_out = 1'b1;
assign local_bb2_var__u58_valid_out = 1'b1;
assign local_bb2_reduction_0_i417_valid_out = 1'b1;
assign local_bb2_var__u52_valid_out = 1'b1;
assign local_bb2__29_i_valid_out = 1'b1;
assign local_bb2__29_i1399_valid_out = 1'b1;
assign local_bb2__29_i851_valid_out = 1'b1;
assign local_bb2__29_i387_valid_out = 1'b1;
assign local_bb2__29_i1307_valid_out = 1'b1;
assign local_bb2__29_i1856_valid_out = 1'b1;
assign local_bb2__29_i759_valid_out = 1'b1;
assign local_bb2__29_i295_valid_out = 1'b1;
assign local_bb2_c0_enter_c0_eni8_stall_in_0 = 1'b0;
assign local_bb2_c0_enter_c0_eni8_stall_in_1 = 1'b0;
assign local_bb2_c0_enter_c0_eni8_stall_in_3 = 1'b0;
assign local_bb2_c0_enter_c0_eni8_stall_in_6 = 1'b0;
assign local_bb2_c0_enter_c0_eni8_stall_in_7 = 1'b0;
assign local_bb2_c0_enter_c0_eni8_stall_in_2 = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_xor_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_xor_i1278_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_xor_i1827_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_xor_i1370_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_xor_i822_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_xor_i266_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_xor_i730_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_xor_i358_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv1_i_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_i1319_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv1_i_i1311_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_i1868_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv1_i_i1860_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_i1411_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv1_i_i1403_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_i863_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv1_i_i855_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_i307_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv1_i_i299_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_i771_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv1_i_i763_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add_i399_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv1_i_i391_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv_i_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv_i_i1402_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv_i_i854_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv_i_i390_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u46_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i1337_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u56_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv_i_i1859_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv_i_i1310_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv_i_i762_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_conv_i_i298_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i1886_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u54_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i1429_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u48_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i881_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u50_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i325_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u60_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i789_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u58_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i417_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u52_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__29_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__29_i1399_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__29_i851_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__29_i387_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__29_i1307_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__29_i1856_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__29_i759_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__29_i295_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_xor_i_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_xor_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_xor_i_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_xor_i1278_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_xor_i1278_consumed_0_NO_SHIFT_REG | ~(local_bb2_xor_i1278_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_xor_i1827_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_xor_i1827_consumed_0_NO_SHIFT_REG | ~(local_bb2_xor_i1827_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_xor_i1370_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_xor_i1370_consumed_0_NO_SHIFT_REG | ~(local_bb2_xor_i1370_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_xor_i822_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_xor_i822_consumed_0_NO_SHIFT_REG | ~(local_bb2_xor_i822_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_xor_i266_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_xor_i266_consumed_0_NO_SHIFT_REG | ~(local_bb2_xor_i266_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_xor_i730_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_xor_i730_consumed_0_NO_SHIFT_REG | ~(local_bb2_xor_i730_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_xor_i358_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_xor_i358_consumed_0_NO_SHIFT_REG | ~(local_bb2_xor_i358_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_add_i_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_add_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_i_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv1_i_i_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv1_i_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv1_i_i_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_add_i1319_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_add_i1319_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_i1319_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv1_i_i1311_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv1_i_i1311_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv1_i_i1311_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_add_i1868_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_add_i1868_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_i1868_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv1_i_i1860_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv1_i_i1860_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv1_i_i1860_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_add_i1411_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_add_i1411_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_i1411_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv1_i_i1403_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv1_i_i1403_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv1_i_i1403_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_add_i863_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_add_i863_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_i863_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv1_i_i855_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv1_i_i855_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv1_i_i855_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_add_i307_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_add_i307_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_i307_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv1_i_i299_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv1_i_i299_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv1_i_i299_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_add_i771_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_add_i771_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_i771_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv1_i_i763_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv1_i_i763_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv1_i_i763_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_add_i399_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_add_i399_consumed_0_NO_SHIFT_REG | ~(local_bb2_add_i399_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv1_i_i391_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv1_i_i391_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv1_i_i391_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv_i_i_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv_i_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv_i_i_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv_i_i1402_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv_i_i1402_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv_i_i1402_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv_i_i854_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv_i_i854_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv_i_i854_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv_i_i390_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv_i_i390_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv_i_i390_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_reduction_0_i_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_reduction_0_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_var__u46_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_var__u46_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u46_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_reduction_0_i1337_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_reduction_0_i1337_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i1337_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_var__u56_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_var__u56_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u56_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv_i_i1859_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv_i_i1859_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv_i_i1859_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv_i_i1310_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv_i_i1310_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv_i_i1310_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv_i_i762_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv_i_i762_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv_i_i762_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_conv_i_i298_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_conv_i_i298_consumed_0_NO_SHIFT_REG | ~(local_bb2_conv_i_i298_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_reduction_0_i1886_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_reduction_0_i1886_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i1886_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_var__u54_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_var__u54_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u54_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_reduction_0_i1429_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_reduction_0_i1429_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i1429_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_var__u48_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_var__u48_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u48_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_reduction_0_i881_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_reduction_0_i881_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i881_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_var__u50_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_var__u50_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u50_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_reduction_0_i325_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_reduction_0_i325_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i325_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_var__u60_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_var__u60_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u60_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_reduction_0_i789_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_reduction_0_i789_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i789_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_var__u58_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_var__u58_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u58_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_reduction_0_i417_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_reduction_0_i417_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i417_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2_var__u52_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2_var__u52_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u52_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2__29_i_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2__29_i_consumed_0_NO_SHIFT_REG | ~(local_bb2__29_i_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2__29_i1399_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2__29_i1399_consumed_0_NO_SHIFT_REG | ~(local_bb2__29_i1399_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2__29_i851_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2__29_i851_consumed_0_NO_SHIFT_REG | ~(local_bb2__29_i851_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2__29_i387_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2__29_i387_consumed_0_NO_SHIFT_REG | ~(local_bb2__29_i387_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2__29_i1307_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2__29_i1307_consumed_0_NO_SHIFT_REG | ~(local_bb2__29_i1307_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2__29_i1856_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2__29_i1856_consumed_0_NO_SHIFT_REG | ~(local_bb2__29_i1856_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2__29_i759_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2__29_i759_consumed_0_NO_SHIFT_REG | ~(local_bb2__29_i759_stall_in)) & local_bb2__29_i387_stall_local);
		local_bb2__29_i295_consumed_0_NO_SHIFT_REG <= (local_bb2__29_i387_inputs_ready & (local_bb2__29_i295_consumed_0_NO_SHIFT_REG | ~(local_bb2__29_i295_stall_in)) & local_bb2__29_i387_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_xor_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_xor_i_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_xor_i_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_xor_i_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_xor_i_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_xor_i_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i),
	.data_out(rnode_166to167_bb2_xor_i_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_xor_i_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_xor_i_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_xor_i_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_xor_i_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_xor_i_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i_stall_in = 1'b0;
assign rnode_166to167_bb2_xor_i_0_NO_SHIFT_REG = rnode_166to167_bb2_xor_i_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_xor_i_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_xor_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_xor_i1278_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1278_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i1278_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1278_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i1278_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1278_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1278_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1278_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_xor_i1278_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_xor_i1278_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_xor_i1278_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_xor_i1278_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_xor_i1278_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i1278),
	.data_out(rnode_166to167_bb2_xor_i1278_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_xor_i1278_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_xor_i1278_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_xor_i1278_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_xor_i1278_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_xor_i1278_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i1278_stall_in = 1'b0;
assign rnode_166to167_bb2_xor_i1278_0_NO_SHIFT_REG = rnode_166to167_bb2_xor_i1278_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_xor_i1278_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_xor_i1278_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_xor_i1827_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1827_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i1827_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1827_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i1827_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1827_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1827_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1827_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_xor_i1827_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_xor_i1827_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_xor_i1827_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_xor_i1827_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_xor_i1827_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i1827),
	.data_out(rnode_166to167_bb2_xor_i1827_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_xor_i1827_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_xor_i1827_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_xor_i1827_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_xor_i1827_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_xor_i1827_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i1827_stall_in = 1'b0;
assign rnode_166to167_bb2_xor_i1827_0_NO_SHIFT_REG = rnode_166to167_bb2_xor_i1827_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_xor_i1827_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_xor_i1827_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_xor_i1370_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1370_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i1370_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1370_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i1370_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1370_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1370_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i1370_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_xor_i1370_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_xor_i1370_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_xor_i1370_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_xor_i1370_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_xor_i1370_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i1370),
	.data_out(rnode_166to167_bb2_xor_i1370_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_xor_i1370_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_xor_i1370_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_xor_i1370_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_xor_i1370_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_xor_i1370_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i1370_stall_in = 1'b0;
assign rnode_166to167_bb2_xor_i1370_0_NO_SHIFT_REG = rnode_166to167_bb2_xor_i1370_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_xor_i1370_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_xor_i1370_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_xor_i822_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i822_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i822_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i822_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i822_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i822_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i822_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i822_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_xor_i822_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_xor_i822_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_xor_i822_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_xor_i822_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_xor_i822_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i822),
	.data_out(rnode_166to167_bb2_xor_i822_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_xor_i822_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_xor_i822_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_xor_i822_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_xor_i822_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_xor_i822_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i822_stall_in = 1'b0;
assign rnode_166to167_bb2_xor_i822_0_NO_SHIFT_REG = rnode_166to167_bb2_xor_i822_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_xor_i822_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_xor_i822_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_xor_i266_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i266_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i266_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i266_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i266_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i266_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i266_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i266_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_xor_i266_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_xor_i266_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_xor_i266_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_xor_i266_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_xor_i266_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i266),
	.data_out(rnode_166to167_bb2_xor_i266_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_xor_i266_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_xor_i266_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_xor_i266_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_xor_i266_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_xor_i266_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i266_stall_in = 1'b0;
assign rnode_166to167_bb2_xor_i266_0_NO_SHIFT_REG = rnode_166to167_bb2_xor_i266_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_xor_i266_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_xor_i266_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_xor_i730_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i730_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i730_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i730_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i730_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i730_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i730_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i730_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_xor_i730_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_xor_i730_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_xor_i730_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_xor_i730_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_xor_i730_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i730),
	.data_out(rnode_166to167_bb2_xor_i730_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_xor_i730_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_xor_i730_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_xor_i730_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_xor_i730_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_xor_i730_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i730_stall_in = 1'b0;
assign rnode_166to167_bb2_xor_i730_0_NO_SHIFT_REG = rnode_166to167_bb2_xor_i730_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_xor_i730_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_xor_i730_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_xor_i358_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i358_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i358_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i358_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_xor_i358_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i358_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i358_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_xor_i358_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_xor_i358_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_xor_i358_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_xor_i358_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_xor_i358_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_xor_i358_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i358),
	.data_out(rnode_166to167_bb2_xor_i358_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_xor_i358_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_xor_i358_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_xor_i358_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_xor_i358_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_xor_i358_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i358_stall_in = 1'b0;
assign rnode_166to167_bb2_xor_i358_0_NO_SHIFT_REG = rnode_166to167_bb2_xor_i358_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_xor_i358_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_xor_i358_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_add_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_add_i_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_add_i_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_add_i_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_add_i_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_add_i_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_add_i),
	.data_out(rnode_166to167_bb2_add_i_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_add_i_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_add_i_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_add_i_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_add_i_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_add_i_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add_i_stall_in = 1'b0;
assign rnode_166to167_bb2_add_i_0_NO_SHIFT_REG = rnode_166to167_bb2_add_i_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_add_i_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_add_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_add_i1319_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1319_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i1319_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1319_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i1319_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1319_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1319_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1319_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_add_i1319_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_add_i1319_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_add_i1319_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_add_i1319_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_add_i1319_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_add_i1319),
	.data_out(rnode_166to167_bb2_add_i1319_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_add_i1319_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_add_i1319_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_add_i1319_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_add_i1319_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_add_i1319_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add_i1319_stall_in = 1'b0;
assign rnode_166to167_bb2_add_i1319_0_NO_SHIFT_REG = rnode_166to167_bb2_add_i1319_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_add_i1319_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_add_i1319_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_add_i1868_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1868_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i1868_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1868_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i1868_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1868_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1868_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1868_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_add_i1868_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_add_i1868_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_add_i1868_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_add_i1868_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_add_i1868_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_add_i1868),
	.data_out(rnode_166to167_bb2_add_i1868_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_add_i1868_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_add_i1868_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_add_i1868_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_add_i1868_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_add_i1868_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add_i1868_stall_in = 1'b0;
assign rnode_166to167_bb2_add_i1868_0_NO_SHIFT_REG = rnode_166to167_bb2_add_i1868_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_add_i1868_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_add_i1868_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_add_i1411_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1411_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i1411_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1411_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i1411_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1411_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1411_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i1411_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_add_i1411_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_add_i1411_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_add_i1411_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_add_i1411_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_add_i1411_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_add_i1411),
	.data_out(rnode_166to167_bb2_add_i1411_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_add_i1411_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_add_i1411_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_add_i1411_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_add_i1411_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_add_i1411_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add_i1411_stall_in = 1'b0;
assign rnode_166to167_bb2_add_i1411_0_NO_SHIFT_REG = rnode_166to167_bb2_add_i1411_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_add_i1411_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_add_i1411_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_add_i863_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i863_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i863_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i863_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i863_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i863_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i863_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i863_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_add_i863_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_add_i863_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_add_i863_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_add_i863_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_add_i863_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_add_i863),
	.data_out(rnode_166to167_bb2_add_i863_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_add_i863_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_add_i863_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_add_i863_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_add_i863_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_add_i863_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add_i863_stall_in = 1'b0;
assign rnode_166to167_bb2_add_i863_0_NO_SHIFT_REG = rnode_166to167_bb2_add_i863_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_add_i863_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_add_i863_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_add_i307_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i307_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i307_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i307_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i307_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i307_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i307_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i307_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_add_i307_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_add_i307_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_add_i307_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_add_i307_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_add_i307_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_add_i307),
	.data_out(rnode_166to167_bb2_add_i307_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_add_i307_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_add_i307_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_add_i307_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_add_i307_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_add_i307_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add_i307_stall_in = 1'b0;
assign rnode_166to167_bb2_add_i307_0_NO_SHIFT_REG = rnode_166to167_bb2_add_i307_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_add_i307_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_add_i307_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_add_i771_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i771_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i771_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i771_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i771_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i771_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i771_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i771_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_add_i771_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_add_i771_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_add_i771_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_add_i771_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_add_i771_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_add_i771),
	.data_out(rnode_166to167_bb2_add_i771_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_add_i771_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_add_i771_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_add_i771_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_add_i771_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_add_i771_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add_i771_stall_in = 1'b0;
assign rnode_166to167_bb2_add_i771_0_NO_SHIFT_REG = rnode_166to167_bb2_add_i771_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_add_i771_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_add_i771_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_add_i399_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i399_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i399_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i399_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_166to167_bb2_add_i399_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i399_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i399_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_add_i399_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_add_i399_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_add_i399_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_add_i399_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_add_i399_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_add_i399_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_add_i399),
	.data_out(rnode_166to167_bb2_add_i399_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_add_i399_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_add_i399_0_reg_167_fifo.DATA_WIDTH = 32;
defparam rnode_166to167_bb2_add_i399_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_add_i399_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_add_i399_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add_i399_stall_in = 1'b0;
assign rnode_166to167_bb2_add_i399_0_NO_SHIFT_REG = rnode_166to167_bb2_add_i399_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_add_i399_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_add_i399_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb2_mul_i_i_inputs_ready;
 reg local_bb2_mul_i_i_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul_i_i_stall_in_0;
 reg local_bb2_mul_i_i_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i_stall_in_1;
wire local_bb2_mul_i_i_output_regs_ready;
wire [63:0] local_bb2_mul_i_i;
 reg local_bb2_mul_i_i_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul_i_i_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i_causedstall;

acl_int_mult64s_s5 int_module_local_bb2_mul_i_i (
	.clock(clock),
	.dataa(local_bb2_conv1_i_i),
	.datab(local_bb2_conv_i_i),
	.enable(local_bb2_mul_i_i_output_regs_ready),
	.result(local_bb2_mul_i_i)
);

defparam int_module_local_bb2_mul_i_i.INPUT1_WIDTH = 24;
defparam int_module_local_bb2_mul_i_i.INPUT2_WIDTH = 24;

assign local_bb2_mul_i_i_inputs_ready = 1'b1;
assign local_bb2_mul_i_i_output_regs_ready = 1'b1;
assign local_bb2_conv1_i_i_stall_in = 1'b0;
assign local_bb2_conv_i_i_stall_in = 1'b0;
assign local_bb2_mul_i_i_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i_output_regs_ready)
		begin
			local_bb2_mul_i_i_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul_i_i_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i_output_regs_ready)
		begin
			local_bb2_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_mul_i_i_stall_in_0))
			begin
				local_bb2_mul_i_i_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul_i_i_stall_in_1))
			begin
				local_bb2_mul_i_i_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul_i_i1404_inputs_ready;
 reg local_bb2_mul_i_i1404_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul_i_i1404_stall_in_0;
 reg local_bb2_mul_i_i1404_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i1404_stall_in_1;
wire local_bb2_mul_i_i1404_output_regs_ready;
wire [63:0] local_bb2_mul_i_i1404;
 reg local_bb2_mul_i_i1404_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul_i_i1404_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i1404_causedstall;

acl_int_mult64s_s5 int_module_local_bb2_mul_i_i1404 (
	.clock(clock),
	.dataa(local_bb2_conv1_i_i1403),
	.datab(local_bb2_conv_i_i1402),
	.enable(local_bb2_mul_i_i1404_output_regs_ready),
	.result(local_bb2_mul_i_i1404)
);

defparam int_module_local_bb2_mul_i_i1404.INPUT1_WIDTH = 24;
defparam int_module_local_bb2_mul_i_i1404.INPUT2_WIDTH = 24;

assign local_bb2_mul_i_i1404_inputs_ready = 1'b1;
assign local_bb2_mul_i_i1404_output_regs_ready = 1'b1;
assign local_bb2_conv1_i_i1403_stall_in = 1'b0;
assign local_bb2_conv_i_i1402_stall_in = 1'b0;
assign local_bb2_mul_i_i1404_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i1404_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i1404_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i1404_output_regs_ready)
		begin
			local_bb2_mul_i_i1404_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i1404_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul_i_i1404_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i1404_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i1404_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i1404_output_regs_ready)
		begin
			local_bb2_mul_i_i1404_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i1404_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_mul_i_i1404_stall_in_0))
			begin
				local_bb2_mul_i_i1404_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul_i_i1404_stall_in_1))
			begin
				local_bb2_mul_i_i1404_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul_i_i856_inputs_ready;
 reg local_bb2_mul_i_i856_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul_i_i856_stall_in_0;
 reg local_bb2_mul_i_i856_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i856_stall_in_1;
wire local_bb2_mul_i_i856_output_regs_ready;
wire [63:0] local_bb2_mul_i_i856;
 reg local_bb2_mul_i_i856_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul_i_i856_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i856_causedstall;

acl_int_mult64s_s5 int_module_local_bb2_mul_i_i856 (
	.clock(clock),
	.dataa(local_bb2_conv1_i_i855),
	.datab(local_bb2_conv_i_i854),
	.enable(local_bb2_mul_i_i856_output_regs_ready),
	.result(local_bb2_mul_i_i856)
);

defparam int_module_local_bb2_mul_i_i856.INPUT1_WIDTH = 24;
defparam int_module_local_bb2_mul_i_i856.INPUT2_WIDTH = 24;

assign local_bb2_mul_i_i856_inputs_ready = 1'b1;
assign local_bb2_mul_i_i856_output_regs_ready = 1'b1;
assign local_bb2_conv1_i_i855_stall_in = 1'b0;
assign local_bb2_conv_i_i854_stall_in = 1'b0;
assign local_bb2_mul_i_i856_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i856_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i856_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i856_output_regs_ready)
		begin
			local_bb2_mul_i_i856_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i856_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul_i_i856_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i856_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i856_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i856_output_regs_ready)
		begin
			local_bb2_mul_i_i856_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i856_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_mul_i_i856_stall_in_0))
			begin
				local_bb2_mul_i_i856_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul_i_i856_stall_in_1))
			begin
				local_bb2_mul_i_i856_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul_i_i392_inputs_ready;
 reg local_bb2_mul_i_i392_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul_i_i392_stall_in_0;
 reg local_bb2_mul_i_i392_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i392_stall_in_1;
wire local_bb2_mul_i_i392_output_regs_ready;
wire [63:0] local_bb2_mul_i_i392;
 reg local_bb2_mul_i_i392_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul_i_i392_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i392_causedstall;

acl_int_mult64s_s5 int_module_local_bb2_mul_i_i392 (
	.clock(clock),
	.dataa(local_bb2_conv1_i_i391),
	.datab(local_bb2_conv_i_i390),
	.enable(local_bb2_mul_i_i392_output_regs_ready),
	.result(local_bb2_mul_i_i392)
);

defparam int_module_local_bb2_mul_i_i392.INPUT1_WIDTH = 24;
defparam int_module_local_bb2_mul_i_i392.INPUT2_WIDTH = 24;

assign local_bb2_mul_i_i392_inputs_ready = 1'b1;
assign local_bb2_mul_i_i392_output_regs_ready = 1'b1;
assign local_bb2_conv1_i_i391_stall_in = 1'b0;
assign local_bb2_conv_i_i390_stall_in = 1'b0;
assign local_bb2_mul_i_i392_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i392_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i392_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i392_output_regs_ready)
		begin
			local_bb2_mul_i_i392_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i392_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul_i_i392_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i392_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i392_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i392_output_regs_ready)
		begin
			local_bb2_mul_i_i392_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i392_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_mul_i_i392_stall_in_0))
			begin
				local_bb2_mul_i_i392_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul_i_i392_stall_in_1))
			begin
				local_bb2_mul_i_i392_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_reduction_0_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_reduction_0_i_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_reduction_0_i_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_reduction_0_i_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_reduction_0_i_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_reduction_0_i_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i),
	.data_out(rnode_166to167_bb2_reduction_0_i_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_reduction_0_i_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_reduction_0_i_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_reduction_0_i_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_reduction_0_i_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_reduction_0_i_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i_stall_in = 1'b0;
assign rnode_166to167_bb2_reduction_0_i_0_NO_SHIFT_REG = rnode_166to167_bb2_reduction_0_i_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_reduction_0_i_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_reduction_0_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_var__u46_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u46_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u46_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u46_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u46_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u46_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u46_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u46_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_var__u46_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_var__u46_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_var__u46_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_var__u46_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_var__u46_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_var__u46),
	.data_out(rnode_166to167_bb2_var__u46_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_var__u46_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_var__u46_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_var__u46_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_var__u46_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_var__u46_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u46_stall_in = 1'b0;
assign rnode_166to167_bb2_var__u46_0_NO_SHIFT_REG = rnode_166to167_bb2_var__u46_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_var__u46_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_var__u46_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_reduction_0_i1337_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1337_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1337_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1337_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1337_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1337_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1337_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1337_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_reduction_0_i1337_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_reduction_0_i1337_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_reduction_0_i1337_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_reduction_0_i1337_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_reduction_0_i1337_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i1337),
	.data_out(rnode_166to167_bb2_reduction_0_i1337_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_reduction_0_i1337_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_reduction_0_i1337_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_reduction_0_i1337_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_reduction_0_i1337_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_reduction_0_i1337_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i1337_stall_in = 1'b0;
assign rnode_166to167_bb2_reduction_0_i1337_0_NO_SHIFT_REG = rnode_166to167_bb2_reduction_0_i1337_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_reduction_0_i1337_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_reduction_0_i1337_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_var__u56_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u56_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u56_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u56_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u56_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u56_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u56_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u56_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_var__u56_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_var__u56_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_var__u56_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_var__u56_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_var__u56_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_var__u56),
	.data_out(rnode_166to167_bb2_var__u56_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_var__u56_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_var__u56_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_var__u56_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_var__u56_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_var__u56_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u56_stall_in = 1'b0;
assign rnode_166to167_bb2_var__u56_0_NO_SHIFT_REG = rnode_166to167_bb2_var__u56_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_var__u56_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_var__u56_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements a registered operation.
// 
wire local_bb2_mul_i_i1861_inputs_ready;
 reg local_bb2_mul_i_i1861_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul_i_i1861_stall_in_0;
 reg local_bb2_mul_i_i1861_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i1861_stall_in_1;
wire local_bb2_mul_i_i1861_output_regs_ready;
wire [63:0] local_bb2_mul_i_i1861;
 reg local_bb2_mul_i_i1861_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul_i_i1861_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i1861_causedstall;

acl_int_mult64s_s5 int_module_local_bb2_mul_i_i1861 (
	.clock(clock),
	.dataa(local_bb2_conv1_i_i1860),
	.datab(local_bb2_conv_i_i1859),
	.enable(local_bb2_mul_i_i1861_output_regs_ready),
	.result(local_bb2_mul_i_i1861)
);

defparam int_module_local_bb2_mul_i_i1861.INPUT1_WIDTH = 24;
defparam int_module_local_bb2_mul_i_i1861.INPUT2_WIDTH = 24;

assign local_bb2_mul_i_i1861_inputs_ready = 1'b1;
assign local_bb2_mul_i_i1861_output_regs_ready = 1'b1;
assign local_bb2_conv1_i_i1860_stall_in = 1'b0;
assign local_bb2_conv_i_i1859_stall_in = 1'b0;
assign local_bb2_mul_i_i1861_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i1861_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i1861_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i1861_output_regs_ready)
		begin
			local_bb2_mul_i_i1861_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i1861_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul_i_i1861_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i1861_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i1861_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i1861_output_regs_ready)
		begin
			local_bb2_mul_i_i1861_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i1861_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_mul_i_i1861_stall_in_0))
			begin
				local_bb2_mul_i_i1861_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul_i_i1861_stall_in_1))
			begin
				local_bb2_mul_i_i1861_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul_i_i1312_inputs_ready;
 reg local_bb2_mul_i_i1312_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul_i_i1312_stall_in_0;
 reg local_bb2_mul_i_i1312_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i1312_stall_in_1;
wire local_bb2_mul_i_i1312_output_regs_ready;
wire [63:0] local_bb2_mul_i_i1312;
 reg local_bb2_mul_i_i1312_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul_i_i1312_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i1312_causedstall;

acl_int_mult64s_s5 int_module_local_bb2_mul_i_i1312 (
	.clock(clock),
	.dataa(local_bb2_conv1_i_i1311),
	.datab(local_bb2_conv_i_i1310),
	.enable(local_bb2_mul_i_i1312_output_regs_ready),
	.result(local_bb2_mul_i_i1312)
);

defparam int_module_local_bb2_mul_i_i1312.INPUT1_WIDTH = 24;
defparam int_module_local_bb2_mul_i_i1312.INPUT2_WIDTH = 24;

assign local_bb2_mul_i_i1312_inputs_ready = 1'b1;
assign local_bb2_mul_i_i1312_output_regs_ready = 1'b1;
assign local_bb2_conv1_i_i1311_stall_in = 1'b0;
assign local_bb2_conv_i_i1310_stall_in = 1'b0;
assign local_bb2_mul_i_i1312_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i1312_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i1312_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i1312_output_regs_ready)
		begin
			local_bb2_mul_i_i1312_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i1312_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul_i_i1312_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i1312_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i1312_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i1312_output_regs_ready)
		begin
			local_bb2_mul_i_i1312_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i1312_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_mul_i_i1312_stall_in_0))
			begin
				local_bb2_mul_i_i1312_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul_i_i1312_stall_in_1))
			begin
				local_bb2_mul_i_i1312_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul_i_i764_inputs_ready;
 reg local_bb2_mul_i_i764_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul_i_i764_stall_in_0;
 reg local_bb2_mul_i_i764_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i764_stall_in_1;
wire local_bb2_mul_i_i764_output_regs_ready;
wire [63:0] local_bb2_mul_i_i764;
 reg local_bb2_mul_i_i764_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul_i_i764_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i764_causedstall;

acl_int_mult64s_s5 int_module_local_bb2_mul_i_i764 (
	.clock(clock),
	.dataa(local_bb2_conv1_i_i763),
	.datab(local_bb2_conv_i_i762),
	.enable(local_bb2_mul_i_i764_output_regs_ready),
	.result(local_bb2_mul_i_i764)
);

defparam int_module_local_bb2_mul_i_i764.INPUT1_WIDTH = 24;
defparam int_module_local_bb2_mul_i_i764.INPUT2_WIDTH = 24;

assign local_bb2_mul_i_i764_inputs_ready = 1'b1;
assign local_bb2_mul_i_i764_output_regs_ready = 1'b1;
assign local_bb2_conv1_i_i763_stall_in = 1'b0;
assign local_bb2_conv_i_i762_stall_in = 1'b0;
assign local_bb2_mul_i_i764_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i764_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i764_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i764_output_regs_ready)
		begin
			local_bb2_mul_i_i764_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i764_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul_i_i764_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i764_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i764_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i764_output_regs_ready)
		begin
			local_bb2_mul_i_i764_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i764_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_mul_i_i764_stall_in_0))
			begin
				local_bb2_mul_i_i764_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul_i_i764_stall_in_1))
			begin
				local_bb2_mul_i_i764_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb2_mul_i_i300_inputs_ready;
 reg local_bb2_mul_i_i300_valid_out_0_NO_SHIFT_REG;
wire local_bb2_mul_i_i300_stall_in_0;
 reg local_bb2_mul_i_i300_valid_out_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i300_stall_in_1;
wire local_bb2_mul_i_i300_output_regs_ready;
wire [63:0] local_bb2_mul_i_i300;
 reg local_bb2_mul_i_i300_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb2_mul_i_i300_valid_pipe_1_NO_SHIFT_REG;
wire local_bb2_mul_i_i300_causedstall;

acl_int_mult64s_s5 int_module_local_bb2_mul_i_i300 (
	.clock(clock),
	.dataa(local_bb2_conv1_i_i299),
	.datab(local_bb2_conv_i_i298),
	.enable(local_bb2_mul_i_i300_output_regs_ready),
	.result(local_bb2_mul_i_i300)
);

defparam int_module_local_bb2_mul_i_i300.INPUT1_WIDTH = 24;
defparam int_module_local_bb2_mul_i_i300.INPUT2_WIDTH = 24;

assign local_bb2_mul_i_i300_inputs_ready = 1'b1;
assign local_bb2_mul_i_i300_output_regs_ready = 1'b1;
assign local_bb2_conv1_i_i299_stall_in = 1'b0;
assign local_bb2_conv_i_i298_stall_in = 1'b0;
assign local_bb2_mul_i_i300_causedstall = (1'b1 && (1'b0 && !(1'b0)));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i300_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i300_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i300_output_regs_ready)
		begin
			local_bb2_mul_i_i300_valid_pipe_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i300_valid_pipe_1_NO_SHIFT_REG <= local_bb2_mul_i_i300_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_mul_i_i300_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_mul_i_i300_valid_out_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_mul_i_i300_output_regs_ready)
		begin
			local_bb2_mul_i_i300_valid_out_0_NO_SHIFT_REG <= 1'b1;
			local_bb2_mul_i_i300_valid_out_1_NO_SHIFT_REG <= 1'b1;
		end
		else
		begin
			if (~(local_bb2_mul_i_i300_stall_in_0))
			begin
				local_bb2_mul_i_i300_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_mul_i_i300_stall_in_1))
			begin
				local_bb2_mul_i_i300_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_reduction_0_i1886_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1886_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1886_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1886_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1886_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1886_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1886_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1886_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_reduction_0_i1886_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_reduction_0_i1886_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_reduction_0_i1886_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_reduction_0_i1886_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_reduction_0_i1886_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i1886),
	.data_out(rnode_166to167_bb2_reduction_0_i1886_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_reduction_0_i1886_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_reduction_0_i1886_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_reduction_0_i1886_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_reduction_0_i1886_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_reduction_0_i1886_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i1886_stall_in = 1'b0;
assign rnode_166to167_bb2_reduction_0_i1886_0_NO_SHIFT_REG = rnode_166to167_bb2_reduction_0_i1886_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_reduction_0_i1886_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_reduction_0_i1886_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_var__u54_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u54_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u54_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u54_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u54_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u54_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u54_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u54_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_var__u54_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_var__u54_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_var__u54_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_var__u54_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_var__u54_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_var__u54),
	.data_out(rnode_166to167_bb2_var__u54_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_var__u54_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_var__u54_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_var__u54_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_var__u54_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_var__u54_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u54_stall_in = 1'b0;
assign rnode_166to167_bb2_var__u54_0_NO_SHIFT_REG = rnode_166to167_bb2_var__u54_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_var__u54_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_var__u54_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_reduction_0_i1429_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1429_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1429_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1429_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1429_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1429_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1429_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i1429_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_reduction_0_i1429_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_reduction_0_i1429_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_reduction_0_i1429_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_reduction_0_i1429_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_reduction_0_i1429_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i1429),
	.data_out(rnode_166to167_bb2_reduction_0_i1429_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_reduction_0_i1429_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_reduction_0_i1429_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_reduction_0_i1429_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_reduction_0_i1429_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_reduction_0_i1429_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i1429_stall_in = 1'b0;
assign rnode_166to167_bb2_reduction_0_i1429_0_NO_SHIFT_REG = rnode_166to167_bb2_reduction_0_i1429_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_reduction_0_i1429_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_reduction_0_i1429_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_var__u48_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u48_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u48_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u48_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u48_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u48_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u48_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u48_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_var__u48_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_var__u48_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_var__u48_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_var__u48_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_var__u48_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_var__u48),
	.data_out(rnode_166to167_bb2_var__u48_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_var__u48_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_var__u48_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_var__u48_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_var__u48_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_var__u48_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u48_stall_in = 1'b0;
assign rnode_166to167_bb2_var__u48_0_NO_SHIFT_REG = rnode_166to167_bb2_var__u48_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_var__u48_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_var__u48_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_reduction_0_i881_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i881_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i881_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i881_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i881_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i881_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i881_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i881_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_reduction_0_i881_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_reduction_0_i881_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_reduction_0_i881_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_reduction_0_i881_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_reduction_0_i881_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i881),
	.data_out(rnode_166to167_bb2_reduction_0_i881_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_reduction_0_i881_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_reduction_0_i881_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_reduction_0_i881_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_reduction_0_i881_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_reduction_0_i881_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i881_stall_in = 1'b0;
assign rnode_166to167_bb2_reduction_0_i881_0_NO_SHIFT_REG = rnode_166to167_bb2_reduction_0_i881_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_reduction_0_i881_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_reduction_0_i881_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_var__u50_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u50_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u50_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u50_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u50_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u50_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u50_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u50_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_var__u50_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_var__u50_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_var__u50_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_var__u50_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_var__u50_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_var__u50),
	.data_out(rnode_166to167_bb2_var__u50_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_var__u50_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_var__u50_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_var__u50_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_var__u50_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_var__u50_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u50_stall_in = 1'b0;
assign rnode_166to167_bb2_var__u50_0_NO_SHIFT_REG = rnode_166to167_bb2_var__u50_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_var__u50_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_var__u50_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_reduction_0_i325_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i325_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i325_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i325_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i325_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i325_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i325_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i325_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_reduction_0_i325_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_reduction_0_i325_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_reduction_0_i325_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_reduction_0_i325_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_reduction_0_i325_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i325),
	.data_out(rnode_166to167_bb2_reduction_0_i325_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_reduction_0_i325_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_reduction_0_i325_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_reduction_0_i325_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_reduction_0_i325_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_reduction_0_i325_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i325_stall_in = 1'b0;
assign rnode_166to167_bb2_reduction_0_i325_0_NO_SHIFT_REG = rnode_166to167_bb2_reduction_0_i325_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_reduction_0_i325_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_reduction_0_i325_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_var__u60_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u60_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u60_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u60_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u60_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u60_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u60_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u60_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_var__u60_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_var__u60_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_var__u60_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_var__u60_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_var__u60_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_var__u60),
	.data_out(rnode_166to167_bb2_var__u60_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_var__u60_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_var__u60_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_var__u60_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_var__u60_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_var__u60_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u60_stall_in = 1'b0;
assign rnode_166to167_bb2_var__u60_0_NO_SHIFT_REG = rnode_166to167_bb2_var__u60_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_var__u60_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_var__u60_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_reduction_0_i789_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i789_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i789_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i789_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i789_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i789_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i789_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i789_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_reduction_0_i789_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_reduction_0_i789_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_reduction_0_i789_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_reduction_0_i789_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_reduction_0_i789_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i789),
	.data_out(rnode_166to167_bb2_reduction_0_i789_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_reduction_0_i789_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_reduction_0_i789_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_reduction_0_i789_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_reduction_0_i789_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_reduction_0_i789_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i789_stall_in = 1'b0;
assign rnode_166to167_bb2_reduction_0_i789_0_NO_SHIFT_REG = rnode_166to167_bb2_reduction_0_i789_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_reduction_0_i789_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_reduction_0_i789_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_var__u58_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u58_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u58_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u58_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u58_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u58_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u58_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u58_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_var__u58_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_var__u58_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_var__u58_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_var__u58_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_var__u58_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_var__u58),
	.data_out(rnode_166to167_bb2_var__u58_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_var__u58_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_var__u58_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_var__u58_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_var__u58_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_var__u58_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u58_stall_in = 1'b0;
assign rnode_166to167_bb2_var__u58_0_NO_SHIFT_REG = rnode_166to167_bb2_var__u58_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_var__u58_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_var__u58_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_reduction_0_i417_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i417_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i417_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i417_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i417_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i417_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i417_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_reduction_0_i417_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_reduction_0_i417_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_reduction_0_i417_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_reduction_0_i417_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_reduction_0_i417_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_reduction_0_i417_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i417),
	.data_out(rnode_166to167_bb2_reduction_0_i417_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_reduction_0_i417_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_reduction_0_i417_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_reduction_0_i417_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_reduction_0_i417_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_reduction_0_i417_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i417_stall_in = 1'b0;
assign rnode_166to167_bb2_reduction_0_i417_0_NO_SHIFT_REG = rnode_166to167_bb2_reduction_0_i417_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_reduction_0_i417_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_reduction_0_i417_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2_var__u52_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u52_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u52_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u52_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u52_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u52_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u52_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2_var__u52_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2_var__u52_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2_var__u52_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2_var__u52_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2_var__u52_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2_var__u52_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2_var__u52),
	.data_out(rnode_166to167_bb2_var__u52_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2_var__u52_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2_var__u52_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2_var__u52_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2_var__u52_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2_var__u52_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u52_stall_in = 1'b0;
assign rnode_166to167_bb2_var__u52_0_NO_SHIFT_REG = rnode_166to167_bb2_var__u52_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2_var__u52_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2_var__u52_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2__29_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2__29_i_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2__29_i_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2__29_i_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2__29_i_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2__29_i_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2__29_i),
	.data_out(rnode_166to167_bb2__29_i_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2__29_i_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2__29_i_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2__29_i_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2__29_i_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2__29_i_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__29_i_stall_in = 1'b0;
assign rnode_166to167_bb2__29_i_0_NO_SHIFT_REG = rnode_166to167_bb2__29_i_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2__29_i_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2__29_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2__29_i1399_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1399_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1399_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1399_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1399_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1399_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1399_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1399_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2__29_i1399_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2__29_i1399_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2__29_i1399_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2__29_i1399_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2__29_i1399_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2__29_i1399),
	.data_out(rnode_166to167_bb2__29_i1399_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2__29_i1399_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2__29_i1399_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2__29_i1399_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2__29_i1399_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2__29_i1399_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__29_i1399_stall_in = 1'b0;
assign rnode_166to167_bb2__29_i1399_0_NO_SHIFT_REG = rnode_166to167_bb2__29_i1399_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2__29_i1399_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2__29_i1399_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2__29_i851_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i851_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i851_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i851_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i851_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i851_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i851_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i851_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2__29_i851_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2__29_i851_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2__29_i851_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2__29_i851_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2__29_i851_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2__29_i851),
	.data_out(rnode_166to167_bb2__29_i851_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2__29_i851_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2__29_i851_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2__29_i851_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2__29_i851_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2__29_i851_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__29_i851_stall_in = 1'b0;
assign rnode_166to167_bb2__29_i851_0_NO_SHIFT_REG = rnode_166to167_bb2__29_i851_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2__29_i851_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2__29_i851_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2__29_i387_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i387_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i387_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i387_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i387_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i387_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i387_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i387_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2__29_i387_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2__29_i387_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2__29_i387_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2__29_i387_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2__29_i387_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2__29_i387),
	.data_out(rnode_166to167_bb2__29_i387_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2__29_i387_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2__29_i387_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2__29_i387_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2__29_i387_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2__29_i387_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__29_i387_stall_in = 1'b0;
assign rnode_166to167_bb2__29_i387_0_NO_SHIFT_REG = rnode_166to167_bb2__29_i387_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2__29_i387_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2__29_i387_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2__29_i1307_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1307_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1307_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1307_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1307_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1307_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1307_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1307_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2__29_i1307_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2__29_i1307_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2__29_i1307_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2__29_i1307_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2__29_i1307_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2__29_i1307),
	.data_out(rnode_166to167_bb2__29_i1307_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2__29_i1307_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2__29_i1307_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2__29_i1307_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2__29_i1307_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2__29_i1307_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__29_i1307_stall_in = 1'b0;
assign rnode_166to167_bb2__29_i1307_0_NO_SHIFT_REG = rnode_166to167_bb2__29_i1307_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2__29_i1307_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2__29_i1307_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2__29_i1856_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1856_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1856_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1856_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1856_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1856_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1856_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i1856_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2__29_i1856_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2__29_i1856_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2__29_i1856_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2__29_i1856_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2__29_i1856_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2__29_i1856),
	.data_out(rnode_166to167_bb2__29_i1856_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2__29_i1856_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2__29_i1856_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2__29_i1856_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2__29_i1856_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2__29_i1856_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__29_i1856_stall_in = 1'b0;
assign rnode_166to167_bb2__29_i1856_0_NO_SHIFT_REG = rnode_166to167_bb2__29_i1856_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2__29_i1856_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2__29_i1856_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2__29_i759_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i759_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i759_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i759_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i759_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i759_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i759_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i759_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2__29_i759_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2__29_i759_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2__29_i759_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2__29_i759_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2__29_i759_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2__29_i759),
	.data_out(rnode_166to167_bb2__29_i759_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2__29_i759_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2__29_i759_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2__29_i759_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2__29_i759_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2__29_i759_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__29_i759_stall_in = 1'b0;
assign rnode_166to167_bb2__29_i759_0_NO_SHIFT_REG = rnode_166to167_bb2__29_i759_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2__29_i759_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2__29_i759_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_166to167_bb2__29_i295_0_valid_out_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i295_0_stall_in_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i295_0_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i295_0_reg_167_inputs_ready_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i295_0_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i295_0_valid_out_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i295_0_stall_in_reg_167_NO_SHIFT_REG;
 logic rnode_166to167_bb2__29_i295_0_stall_out_reg_167_NO_SHIFT_REG;

acl_data_fifo rnode_166to167_bb2__29_i295_0_reg_167_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_166to167_bb2__29_i295_0_reg_167_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_166to167_bb2__29_i295_0_stall_in_reg_167_NO_SHIFT_REG),
	.valid_out(rnode_166to167_bb2__29_i295_0_valid_out_reg_167_NO_SHIFT_REG),
	.stall_out(rnode_166to167_bb2__29_i295_0_stall_out_reg_167_NO_SHIFT_REG),
	.data_in(local_bb2__29_i295),
	.data_out(rnode_166to167_bb2__29_i295_0_reg_167_NO_SHIFT_REG)
);

defparam rnode_166to167_bb2__29_i295_0_reg_167_fifo.DEPTH = 1;
defparam rnode_166to167_bb2__29_i295_0_reg_167_fifo.DATA_WIDTH = 1;
defparam rnode_166to167_bb2__29_i295_0_reg_167_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_166to167_bb2__29_i295_0_reg_167_fifo.IMPL = "shift_reg";

assign rnode_166to167_bb2__29_i295_0_reg_167_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__29_i295_stall_in = 1'b0;
assign rnode_166to167_bb2__29_i295_0_NO_SHIFT_REG = rnode_166to167_bb2__29_i295_0_reg_167_NO_SHIFT_REG;
assign rnode_166to167_bb2__29_i295_0_stall_in_reg_167_NO_SHIFT_REG = 1'b0;
assign rnode_166to167_bb2__29_i295_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_xor_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_xor_i_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_xor_i_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_xor_i_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_xor_i_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_xor_i_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_xor_i_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_xor_i_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_xor_i_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_xor_i_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_167to169_bb2_xor_i_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_xor_i_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_xor_i_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_xor_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i_0_NO_SHIFT_REG = rnode_167to169_bb2_xor_i_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_xor_i_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_xor_i1278_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1278_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i1278_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1278_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i1278_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1278_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1278_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1278_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_xor_i1278_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_xor_i1278_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_xor_i1278_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_xor_i1278_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_xor_i1278_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_xor_i1278_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_xor_i1278_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_xor_i1278_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_xor_i1278_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_167to169_bb2_xor_i1278_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_xor_i1278_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_xor_i1278_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_xor_i1278_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i1278_0_NO_SHIFT_REG = rnode_167to169_bb2_xor_i1278_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_xor_i1278_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i1278_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_xor_i1827_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1827_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i1827_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1827_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i1827_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1827_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1827_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1827_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_xor_i1827_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_xor_i1827_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_xor_i1827_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_xor_i1827_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_xor_i1827_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_xor_i1827_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_xor_i1827_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_xor_i1827_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_xor_i1827_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_167to169_bb2_xor_i1827_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_xor_i1827_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_xor_i1827_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_xor_i1827_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i1827_0_NO_SHIFT_REG = rnode_167to169_bb2_xor_i1827_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_xor_i1827_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i1827_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_xor_i1370_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1370_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i1370_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1370_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i1370_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1370_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1370_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i1370_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_xor_i1370_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_xor_i1370_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_xor_i1370_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_xor_i1370_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_xor_i1370_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_xor_i1370_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_xor_i1370_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_xor_i1370_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_xor_i1370_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_167to169_bb2_xor_i1370_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_xor_i1370_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_xor_i1370_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_xor_i1370_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i1370_0_NO_SHIFT_REG = rnode_167to169_bb2_xor_i1370_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_xor_i1370_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i1370_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_xor_i822_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i822_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i822_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i822_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i822_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i822_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i822_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i822_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_xor_i822_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_xor_i822_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_xor_i822_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_xor_i822_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_xor_i822_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_xor_i822_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_xor_i822_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_xor_i822_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_xor_i822_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_167to169_bb2_xor_i822_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_xor_i822_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_xor_i822_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_xor_i822_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i822_0_NO_SHIFT_REG = rnode_167to169_bb2_xor_i822_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_xor_i822_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i822_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_xor_i266_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i266_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i266_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i266_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i266_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i266_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i266_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i266_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_xor_i266_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_xor_i266_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_xor_i266_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_xor_i266_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_xor_i266_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_xor_i266_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_xor_i266_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_xor_i266_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_xor_i266_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_167to169_bb2_xor_i266_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_xor_i266_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_xor_i266_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_xor_i266_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i266_0_NO_SHIFT_REG = rnode_167to169_bb2_xor_i266_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_xor_i266_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i266_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_xor_i730_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i730_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i730_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i730_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i730_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i730_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i730_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i730_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_xor_i730_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_xor_i730_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_xor_i730_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_xor_i730_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_xor_i730_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_xor_i730_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_xor_i730_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_xor_i730_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_xor_i730_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_167to169_bb2_xor_i730_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_xor_i730_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_xor_i730_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_xor_i730_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i730_0_NO_SHIFT_REG = rnode_167to169_bb2_xor_i730_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_xor_i730_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i730_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_xor_i358_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i358_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i358_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i358_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to169_bb2_xor_i358_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i358_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i358_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_xor_i358_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_xor_i358_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_xor_i358_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_xor_i358_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_xor_i358_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_xor_i358_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_xor_i358_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_xor_i358_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_xor_i358_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_xor_i358_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_167to169_bb2_xor_i358_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_xor_i358_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_xor_i358_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_xor_i358_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i358_0_NO_SHIFT_REG = rnode_167to169_bb2_xor_i358_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_xor_i358_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_xor_i358_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_add_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_add_i_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_add_i_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_add_i_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_add_i_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_add_i_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_add_i_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_add_i_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_add_i_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_add_i_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_167to168_bb2_add_i_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_add_i_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_add_i_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_add_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i_0_NO_SHIFT_REG = rnode_167to168_bb2_add_i_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_add_i_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_add_i1319_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1319_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i1319_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1319_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i1319_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1319_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1319_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1319_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_add_i1319_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_add_i1319_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_add_i1319_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_add_i1319_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_add_i1319_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_add_i1319_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_add_i1319_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_add_i1319_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_add_i1319_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_167to168_bb2_add_i1319_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_add_i1319_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_add_i1319_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_add_i1319_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i1319_0_NO_SHIFT_REG = rnode_167to168_bb2_add_i1319_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_add_i1319_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i1319_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_add_i1868_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1868_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i1868_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1868_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i1868_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1868_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1868_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1868_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_add_i1868_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_add_i1868_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_add_i1868_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_add_i1868_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_add_i1868_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_add_i1868_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_add_i1868_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_add_i1868_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_add_i1868_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_167to168_bb2_add_i1868_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_add_i1868_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_add_i1868_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_add_i1868_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i1868_0_NO_SHIFT_REG = rnode_167to168_bb2_add_i1868_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_add_i1868_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i1868_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_add_i1411_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1411_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i1411_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1411_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i1411_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1411_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1411_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i1411_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_add_i1411_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_add_i1411_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_add_i1411_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_add_i1411_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_add_i1411_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_add_i1411_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_add_i1411_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_add_i1411_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_add_i1411_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_167to168_bb2_add_i1411_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_add_i1411_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_add_i1411_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_add_i1411_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i1411_0_NO_SHIFT_REG = rnode_167to168_bb2_add_i1411_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_add_i1411_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i1411_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_add_i863_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i863_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i863_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i863_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i863_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i863_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i863_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i863_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_add_i863_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_add_i863_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_add_i863_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_add_i863_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_add_i863_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_add_i863_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_add_i863_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_add_i863_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_add_i863_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_167to168_bb2_add_i863_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_add_i863_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_add_i863_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_add_i863_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i863_0_NO_SHIFT_REG = rnode_167to168_bb2_add_i863_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_add_i863_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i863_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_add_i307_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i307_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i307_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i307_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i307_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i307_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i307_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i307_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_add_i307_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_add_i307_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_add_i307_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_add_i307_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_add_i307_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_add_i307_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_add_i307_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_add_i307_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_add_i307_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_167to168_bb2_add_i307_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_add_i307_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_add_i307_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_add_i307_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i307_0_NO_SHIFT_REG = rnode_167to168_bb2_add_i307_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_add_i307_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i307_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_add_i771_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i771_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i771_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i771_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i771_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i771_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i771_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i771_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_add_i771_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_add_i771_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_add_i771_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_add_i771_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_add_i771_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_add_i771_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_add_i771_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_add_i771_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_add_i771_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_167to168_bb2_add_i771_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_add_i771_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_add_i771_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_add_i771_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i771_0_NO_SHIFT_REG = rnode_167to168_bb2_add_i771_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_add_i771_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i771_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_add_i399_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i399_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i399_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i399_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_167to168_bb2_add_i399_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i399_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i399_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_add_i399_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_add_i399_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_add_i399_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_add_i399_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_add_i399_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_add_i399_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_add_i399_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_add_i399_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_add_i399_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_add_i399_0_reg_168_fifo.DATA_WIDTH = 32;
defparam rnode_167to168_bb2_add_i399_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_add_i399_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_add_i399_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_add_i399_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i399_0_NO_SHIFT_REG = rnode_167to168_bb2_add_i399_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_add_i399_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_add_i399_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_conv3_i_i_stall_local;
wire [31:0] local_bb2_conv3_i_i;

assign local_bb2_conv3_i_i = local_bb2_mul_i_i[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u62_stall_local;
wire [63:0] local_bb2_var__u62;

assign local_bb2_var__u62 = (local_bb2_mul_i_i >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_conv3_i_i1405_stall_local;
wire [31:0] local_bb2_conv3_i_i1405;

assign local_bb2_conv3_i_i1405 = local_bb2_mul_i_i1404[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u63_stall_local;
wire [63:0] local_bb2_var__u63;

assign local_bb2_var__u63 = (local_bb2_mul_i_i1404 >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_conv3_i_i857_stall_local;
wire [31:0] local_bb2_conv3_i_i857;

assign local_bb2_conv3_i_i857 = local_bb2_mul_i_i856[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u64_stall_local;
wire [63:0] local_bb2_var__u64;

assign local_bb2_var__u64 = (local_bb2_mul_i_i856 >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_conv3_i_i393_stall_local;
wire [31:0] local_bb2_conv3_i_i393;

assign local_bb2_conv3_i_i393 = local_bb2_mul_i_i392[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u65_stall_local;
wire [63:0] local_bb2_var__u65;

assign local_bb2_var__u65 = (local_bb2_mul_i_i392 >> 64'h18);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_reduction_0_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_reduction_0_i_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_reduction_0_i_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_reduction_0_i_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_reduction_0_i_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_reduction_0_i_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_reduction_0_i_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_reduction_0_i_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_reduction_0_i_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_reduction_0_i_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_reduction_0_i_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_reduction_0_i_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_reduction_0_i_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_reduction_0_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i_0_NO_SHIFT_REG = rnode_167to169_bb2_reduction_0_i_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_reduction_0_i_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_var__u46_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u46_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u46_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u46_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u46_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u46_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u46_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u46_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_var__u46_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_var__u46_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_var__u46_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_var__u46_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_var__u46_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_var__u46_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_var__u46_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_var__u46_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_var__u46_0_reg_168_fifo.DATA_WIDTH = 1;
defparam rnode_167to168_bb2_var__u46_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_var__u46_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_var__u46_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_var__u46_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_var__u46_0_NO_SHIFT_REG = rnode_167to168_bb2_var__u46_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_var__u46_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_var__u46_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_reduction_0_i1337_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1337_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1337_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1337_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1337_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1337_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1337_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1337_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_reduction_0_i1337_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_reduction_0_i1337_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_reduction_0_i1337_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_reduction_0_i1337_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_reduction_0_i1337_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_reduction_0_i1337_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_reduction_0_i1337_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_reduction_0_i1337_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_reduction_0_i1337_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_reduction_0_i1337_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_reduction_0_i1337_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_reduction_0_i1337_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_reduction_0_i1337_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i1337_0_NO_SHIFT_REG = rnode_167to169_bb2_reduction_0_i1337_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_reduction_0_i1337_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i1337_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_var__u56_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u56_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u56_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u56_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u56_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u56_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u56_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u56_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_var__u56_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_var__u56_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_var__u56_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_var__u56_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_var__u56_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_var__u56_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_var__u56_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_var__u56_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_var__u56_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_var__u56_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_var__u56_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_var__u56_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_var__u56_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u56_0_NO_SHIFT_REG = rnode_167to169_bb2_var__u56_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_var__u56_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u56_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_conv3_i_i1862_stall_local;
wire [31:0] local_bb2_conv3_i_i1862;

assign local_bb2_conv3_i_i1862 = local_bb2_mul_i_i1861[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u66_stall_local;
wire [63:0] local_bb2_var__u66;

assign local_bb2_var__u66 = (local_bb2_mul_i_i1861 >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_conv3_i_i1313_stall_local;
wire [31:0] local_bb2_conv3_i_i1313;

assign local_bb2_conv3_i_i1313 = local_bb2_mul_i_i1312[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u67_stall_local;
wire [63:0] local_bb2_var__u67;

assign local_bb2_var__u67 = (local_bb2_mul_i_i1312 >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_conv3_i_i765_stall_local;
wire [31:0] local_bb2_conv3_i_i765;

assign local_bb2_conv3_i_i765 = local_bb2_mul_i_i764[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u68_stall_local;
wire [63:0] local_bb2_var__u68;

assign local_bb2_var__u68 = (local_bb2_mul_i_i764 >> 64'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_conv3_i_i301_stall_local;
wire [31:0] local_bb2_conv3_i_i301;

assign local_bb2_conv3_i_i301 = local_bb2_mul_i_i300[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_var__u69_stall_local;
wire [63:0] local_bb2_var__u69;

assign local_bb2_var__u69 = (local_bb2_mul_i_i300 >> 64'h18);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_reduction_0_i1886_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1886_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1886_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1886_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1886_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1886_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1886_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1886_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_reduction_0_i1886_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_reduction_0_i1886_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_reduction_0_i1886_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_reduction_0_i1886_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_reduction_0_i1886_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_reduction_0_i1886_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_reduction_0_i1886_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_reduction_0_i1886_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_reduction_0_i1886_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_reduction_0_i1886_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_reduction_0_i1886_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_reduction_0_i1886_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_reduction_0_i1886_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i1886_0_NO_SHIFT_REG = rnode_167to169_bb2_reduction_0_i1886_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_reduction_0_i1886_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i1886_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_var__u54_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u54_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u54_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u54_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u54_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u54_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u54_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u54_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_var__u54_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_var__u54_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_var__u54_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_var__u54_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_var__u54_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_var__u54_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_var__u54_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_var__u54_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_var__u54_0_reg_168_fifo.DATA_WIDTH = 1;
defparam rnode_167to168_bb2_var__u54_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_var__u54_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_var__u54_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_var__u54_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_var__u54_0_NO_SHIFT_REG = rnode_167to168_bb2_var__u54_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_var__u54_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_var__u54_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_reduction_0_i1429_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1429_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1429_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1429_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1429_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1429_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1429_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i1429_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_reduction_0_i1429_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_reduction_0_i1429_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_reduction_0_i1429_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_reduction_0_i1429_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_reduction_0_i1429_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_reduction_0_i1429_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_reduction_0_i1429_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_reduction_0_i1429_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_reduction_0_i1429_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_reduction_0_i1429_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_reduction_0_i1429_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_reduction_0_i1429_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_reduction_0_i1429_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i1429_0_NO_SHIFT_REG = rnode_167to169_bb2_reduction_0_i1429_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_reduction_0_i1429_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i1429_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_var__u48_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u48_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u48_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u48_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u48_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u48_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u48_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u48_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_var__u48_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_var__u48_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_var__u48_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_var__u48_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_var__u48_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_var__u48_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_var__u48_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_var__u48_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_var__u48_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_var__u48_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_var__u48_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_var__u48_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_var__u48_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u48_0_NO_SHIFT_REG = rnode_167to169_bb2_var__u48_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_var__u48_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u48_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_reduction_0_i881_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i881_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i881_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i881_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i881_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i881_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i881_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i881_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_reduction_0_i881_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_reduction_0_i881_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_reduction_0_i881_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_reduction_0_i881_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_reduction_0_i881_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_reduction_0_i881_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_reduction_0_i881_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_reduction_0_i881_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_reduction_0_i881_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_reduction_0_i881_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_reduction_0_i881_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_reduction_0_i881_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_reduction_0_i881_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i881_0_NO_SHIFT_REG = rnode_167to169_bb2_reduction_0_i881_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_reduction_0_i881_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i881_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_var__u50_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u50_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u50_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u50_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u50_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u50_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u50_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u50_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_var__u50_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_var__u50_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_var__u50_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_var__u50_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_var__u50_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_var__u50_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_var__u50_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_var__u50_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_var__u50_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_var__u50_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_var__u50_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_var__u50_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_var__u50_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u50_0_NO_SHIFT_REG = rnode_167to169_bb2_var__u50_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_var__u50_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u50_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_reduction_0_i325_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i325_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i325_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i325_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i325_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i325_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i325_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i325_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_reduction_0_i325_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_reduction_0_i325_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_reduction_0_i325_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_reduction_0_i325_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_reduction_0_i325_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_reduction_0_i325_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_reduction_0_i325_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_reduction_0_i325_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_reduction_0_i325_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_reduction_0_i325_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_reduction_0_i325_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_reduction_0_i325_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_reduction_0_i325_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i325_0_NO_SHIFT_REG = rnode_167to169_bb2_reduction_0_i325_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_reduction_0_i325_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i325_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_var__u60_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u60_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u60_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u60_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u60_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u60_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u60_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u60_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_var__u60_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_var__u60_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_var__u60_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_var__u60_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_var__u60_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_var__u60_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_var__u60_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_var__u60_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_var__u60_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_var__u60_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_var__u60_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_var__u60_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_var__u60_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u60_0_NO_SHIFT_REG = rnode_167to169_bb2_var__u60_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_var__u60_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u60_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_reduction_0_i789_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i789_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i789_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i789_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i789_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i789_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i789_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i789_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_reduction_0_i789_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_reduction_0_i789_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_reduction_0_i789_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_reduction_0_i789_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_reduction_0_i789_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_reduction_0_i789_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_reduction_0_i789_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_reduction_0_i789_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_reduction_0_i789_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_reduction_0_i789_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_reduction_0_i789_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_reduction_0_i789_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_reduction_0_i789_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i789_0_NO_SHIFT_REG = rnode_167to169_bb2_reduction_0_i789_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_reduction_0_i789_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i789_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_167to168_bb2_var__u58_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u58_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u58_0_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u58_0_reg_168_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u58_0_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u58_0_valid_out_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u58_0_stall_in_reg_168_NO_SHIFT_REG;
 logic rnode_167to168_bb2_var__u58_0_stall_out_reg_168_NO_SHIFT_REG;

acl_data_fifo rnode_167to168_bb2_var__u58_0_reg_168_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to168_bb2_var__u58_0_reg_168_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to168_bb2_var__u58_0_stall_in_reg_168_NO_SHIFT_REG),
	.valid_out(rnode_167to168_bb2_var__u58_0_valid_out_reg_168_NO_SHIFT_REG),
	.stall_out(rnode_167to168_bb2_var__u58_0_stall_out_reg_168_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_var__u58_0_NO_SHIFT_REG),
	.data_out(rnode_167to168_bb2_var__u58_0_reg_168_NO_SHIFT_REG)
);

defparam rnode_167to168_bb2_var__u58_0_reg_168_fifo.DEPTH = 1;
defparam rnode_167to168_bb2_var__u58_0_reg_168_fifo.DATA_WIDTH = 1;
defparam rnode_167to168_bb2_var__u58_0_reg_168_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to168_bb2_var__u58_0_reg_168_fifo.IMPL = "shift_reg";

assign rnode_167to168_bb2_var__u58_0_reg_168_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_var__u58_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_var__u58_0_NO_SHIFT_REG = rnode_167to168_bb2_var__u58_0_reg_168_NO_SHIFT_REG;
assign rnode_167to168_bb2_var__u58_0_stall_in_reg_168_NO_SHIFT_REG = 1'b0;
assign rnode_167to168_bb2_var__u58_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_reduction_0_i417_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i417_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i417_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i417_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i417_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i417_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i417_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_reduction_0_i417_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_reduction_0_i417_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_reduction_0_i417_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_reduction_0_i417_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_reduction_0_i417_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_reduction_0_i417_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_reduction_0_i417_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_reduction_0_i417_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_reduction_0_i417_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_reduction_0_i417_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_reduction_0_i417_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_reduction_0_i417_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_reduction_0_i417_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_reduction_0_i417_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i417_0_NO_SHIFT_REG = rnode_167to169_bb2_reduction_0_i417_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_reduction_0_i417_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_reduction_0_i417_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2_var__u52_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u52_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u52_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u52_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u52_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u52_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u52_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2_var__u52_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2_var__u52_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2_var__u52_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2_var__u52_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2_var__u52_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2_var__u52_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2_var__u52_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2_var__u52_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2_var__u52_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2_var__u52_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2_var__u52_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2_var__u52_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2_var__u52_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2_var__u52_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u52_0_NO_SHIFT_REG = rnode_167to169_bb2_var__u52_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2_var__u52_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2_var__u52_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2__29_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2__29_i_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2__29_i_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2__29_i_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2__29_i_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2__29_i_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2__29_i_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2__29_i_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2__29_i_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2__29_i_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2__29_i_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2__29_i_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2__29_i_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2__29_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i_0_NO_SHIFT_REG = rnode_167to169_bb2__29_i_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2__29_i_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2__29_i1399_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1399_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1399_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1399_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1399_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1399_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1399_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1399_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2__29_i1399_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2__29_i1399_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2__29_i1399_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2__29_i1399_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2__29_i1399_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2__29_i1399_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2__29_i1399_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2__29_i1399_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2__29_i1399_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2__29_i1399_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2__29_i1399_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2__29_i1399_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2__29_i1399_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i1399_0_NO_SHIFT_REG = rnode_167to169_bb2__29_i1399_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2__29_i1399_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i1399_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2__29_i851_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i851_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i851_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i851_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i851_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i851_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i851_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i851_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2__29_i851_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2__29_i851_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2__29_i851_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2__29_i851_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2__29_i851_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2__29_i851_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2__29_i851_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2__29_i851_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2__29_i851_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2__29_i851_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2__29_i851_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2__29_i851_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2__29_i851_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i851_0_NO_SHIFT_REG = rnode_167to169_bb2__29_i851_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2__29_i851_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i851_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2__29_i387_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i387_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i387_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i387_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i387_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i387_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i387_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i387_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2__29_i387_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2__29_i387_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2__29_i387_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2__29_i387_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2__29_i387_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2__29_i387_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2__29_i387_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2__29_i387_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2__29_i387_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2__29_i387_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2__29_i387_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2__29_i387_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2__29_i387_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i387_0_NO_SHIFT_REG = rnode_167to169_bb2__29_i387_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2__29_i387_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i387_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2__29_i1307_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1307_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1307_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1307_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1307_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1307_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1307_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1307_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2__29_i1307_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2__29_i1307_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2__29_i1307_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2__29_i1307_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2__29_i1307_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2__29_i1307_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2__29_i1307_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2__29_i1307_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2__29_i1307_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2__29_i1307_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2__29_i1307_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2__29_i1307_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2__29_i1307_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i1307_0_NO_SHIFT_REG = rnode_167to169_bb2__29_i1307_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2__29_i1307_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i1307_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2__29_i1856_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1856_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1856_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1856_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1856_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1856_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1856_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i1856_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2__29_i1856_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2__29_i1856_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2__29_i1856_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2__29_i1856_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2__29_i1856_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2__29_i1856_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2__29_i1856_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2__29_i1856_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2__29_i1856_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2__29_i1856_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2__29_i1856_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2__29_i1856_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2__29_i1856_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i1856_0_NO_SHIFT_REG = rnode_167to169_bb2__29_i1856_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2__29_i1856_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i1856_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2__29_i759_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i759_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i759_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i759_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i759_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i759_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i759_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i759_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2__29_i759_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2__29_i759_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2__29_i759_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2__29_i759_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2__29_i759_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2__29_i759_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2__29_i759_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2__29_i759_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2__29_i759_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2__29_i759_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2__29_i759_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2__29_i759_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2__29_i759_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i759_0_NO_SHIFT_REG = rnode_167to169_bb2__29_i759_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2__29_i759_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i759_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_167to169_bb2__29_i295_0_valid_out_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i295_0_stall_in_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i295_0_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i295_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i295_0_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i295_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i295_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_167to169_bb2__29_i295_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_167to169_bb2__29_i295_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_167to169_bb2__29_i295_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_167to169_bb2__29_i295_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_167to169_bb2__29_i295_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_167to169_bb2__29_i295_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_166to167_bb2__29_i295_0_NO_SHIFT_REG),
	.data_out(rnode_167to169_bb2__29_i295_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_167to169_bb2__29_i295_0_reg_169_fifo.DEPTH = 2;
defparam rnode_167to169_bb2__29_i295_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_167to169_bb2__29_i295_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_167to169_bb2__29_i295_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_167to169_bb2__29_i295_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_166to167_bb2__29_i295_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i295_0_NO_SHIFT_REG = rnode_167to169_bb2__29_i295_0_reg_169_NO_SHIFT_REG;
assign rnode_167to169_bb2__29_i295_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_167to169_bb2__29_i295_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_xor_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_xor_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_xor_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_xor_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_xor_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_xor_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_xor_i_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_xor_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_xor_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_xor_i_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_xor_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_xor_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_xor_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_xor_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i_0_NO_SHIFT_REG = rnode_169to170_bb2_xor_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_xor_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_xor_i1278_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1278_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i1278_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1278_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i1278_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1278_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1278_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1278_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_xor_i1278_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_xor_i1278_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_xor_i1278_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_xor_i1278_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_xor_i1278_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_xor_i1278_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_xor_i1278_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_xor_i1278_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_xor_i1278_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_xor_i1278_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_xor_i1278_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_xor_i1278_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_xor_i1278_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i1278_0_NO_SHIFT_REG = rnode_169to170_bb2_xor_i1278_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_xor_i1278_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i1278_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_xor_i1827_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1827_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i1827_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1827_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i1827_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1827_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1827_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1827_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_xor_i1827_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_xor_i1827_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_xor_i1827_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_xor_i1827_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_xor_i1827_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_xor_i1827_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_xor_i1827_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_xor_i1827_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_xor_i1827_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_xor_i1827_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_xor_i1827_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_xor_i1827_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_xor_i1827_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i1827_0_NO_SHIFT_REG = rnode_169to170_bb2_xor_i1827_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_xor_i1827_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i1827_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_xor_i1370_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1370_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i1370_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1370_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i1370_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1370_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1370_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i1370_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_xor_i1370_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_xor_i1370_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_xor_i1370_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_xor_i1370_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_xor_i1370_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_xor_i1370_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_xor_i1370_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_xor_i1370_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_xor_i1370_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_xor_i1370_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_xor_i1370_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_xor_i1370_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_xor_i1370_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i1370_0_NO_SHIFT_REG = rnode_169to170_bb2_xor_i1370_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_xor_i1370_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i1370_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_xor_i822_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i822_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i822_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i822_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i822_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i822_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i822_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i822_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_xor_i822_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_xor_i822_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_xor_i822_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_xor_i822_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_xor_i822_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_xor_i822_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_xor_i822_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_xor_i822_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_xor_i822_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_xor_i822_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_xor_i822_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_xor_i822_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_xor_i822_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i822_0_NO_SHIFT_REG = rnode_169to170_bb2_xor_i822_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_xor_i822_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i822_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_xor_i266_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i266_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i266_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i266_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i266_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i266_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i266_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i266_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_xor_i266_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_xor_i266_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_xor_i266_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_xor_i266_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_xor_i266_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_xor_i266_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_xor_i266_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_xor_i266_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_xor_i266_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_xor_i266_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_xor_i266_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_xor_i266_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_xor_i266_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i266_0_NO_SHIFT_REG = rnode_169to170_bb2_xor_i266_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_xor_i266_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i266_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_xor_i730_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i730_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i730_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i730_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i730_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i730_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i730_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i730_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_xor_i730_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_xor_i730_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_xor_i730_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_xor_i730_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_xor_i730_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_xor_i730_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_xor_i730_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_xor_i730_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_xor_i730_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_xor_i730_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_xor_i730_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_xor_i730_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_xor_i730_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i730_0_NO_SHIFT_REG = rnode_169to170_bb2_xor_i730_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_xor_i730_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i730_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_xor_i358_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i358_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i358_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i358_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_xor_i358_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i358_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i358_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_xor_i358_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_xor_i358_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_xor_i358_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_xor_i358_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_xor_i358_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_xor_i358_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_xor_i358_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_xor_i358_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_xor_i358_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_xor_i358_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_xor_i358_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_xor_i358_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_xor_i358_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_xor_i358_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i358_0_NO_SHIFT_REG = rnode_169to170_bb2_xor_i358_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_xor_i358_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_xor_i358_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_add_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_add_i_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_add_i_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_add_i_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_add_i_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_add_i_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_add_i_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_add_i_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_add_i_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_add_i_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_168to169_bb2_add_i_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_add_i_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_add_i_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_add_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i_0_stall_in_0_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i_0_NO_SHIFT_REG = rnode_168to169_bb2_add_i_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i_1_NO_SHIFT_REG = rnode_168to169_bb2_add_i_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i_2_NO_SHIFT_REG = rnode_168to169_bb2_add_i_0_reg_169_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_add_i1319_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1319_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1319_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1319_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1319_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1319_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_add_i1319_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_add_i1319_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_add_i1319_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_add_i1319_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_add_i1319_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_add_i1319_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_add_i1319_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_add_i1319_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_add_i1319_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_168to169_bb2_add_i1319_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_add_i1319_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_add_i1319_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_add_i1319_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1319_0_stall_in_0_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1319_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1319_0_NO_SHIFT_REG = rnode_168to169_bb2_add_i1319_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i1319_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1319_1_NO_SHIFT_REG = rnode_168to169_bb2_add_i1319_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i1319_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1319_2_NO_SHIFT_REG = rnode_168to169_bb2_add_i1319_0_reg_169_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_add_i1868_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1868_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1868_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1868_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1868_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1868_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_add_i1868_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_add_i1868_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_add_i1868_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_add_i1868_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_add_i1868_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_add_i1868_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_add_i1868_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_add_i1868_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_add_i1868_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_168to169_bb2_add_i1868_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_add_i1868_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_add_i1868_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_add_i1868_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1868_0_stall_in_0_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1868_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1868_0_NO_SHIFT_REG = rnode_168to169_bb2_add_i1868_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i1868_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1868_1_NO_SHIFT_REG = rnode_168to169_bb2_add_i1868_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i1868_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1868_2_NO_SHIFT_REG = rnode_168to169_bb2_add_i1868_0_reg_169_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_add_i1411_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1411_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1411_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1411_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i1411_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i1411_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_add_i1411_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_add_i1411_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_add_i1411_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_add_i1411_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_add_i1411_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_add_i1411_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_add_i1411_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_add_i1411_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_add_i1411_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_168to169_bb2_add_i1411_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_add_i1411_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_add_i1411_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_add_i1411_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1411_0_stall_in_0_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1411_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1411_0_NO_SHIFT_REG = rnode_168to169_bb2_add_i1411_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i1411_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1411_1_NO_SHIFT_REG = rnode_168to169_bb2_add_i1411_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i1411_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i1411_2_NO_SHIFT_REG = rnode_168to169_bb2_add_i1411_0_reg_169_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_add_i863_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i863_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i863_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i863_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i863_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i863_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_add_i863_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_add_i863_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_add_i863_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_add_i863_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_add_i863_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_add_i863_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_add_i863_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_add_i863_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_add_i863_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_168to169_bb2_add_i863_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_add_i863_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_add_i863_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_add_i863_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i863_0_stall_in_0_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i863_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i863_0_NO_SHIFT_REG = rnode_168to169_bb2_add_i863_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i863_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i863_1_NO_SHIFT_REG = rnode_168to169_bb2_add_i863_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i863_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i863_2_NO_SHIFT_REG = rnode_168to169_bb2_add_i863_0_reg_169_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_add_i307_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i307_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i307_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i307_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i307_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i307_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_add_i307_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_add_i307_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_add_i307_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_add_i307_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_add_i307_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_add_i307_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_add_i307_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_add_i307_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_add_i307_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_168to169_bb2_add_i307_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_add_i307_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_add_i307_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_add_i307_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i307_0_stall_in_0_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i307_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i307_0_NO_SHIFT_REG = rnode_168to169_bb2_add_i307_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i307_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i307_1_NO_SHIFT_REG = rnode_168to169_bb2_add_i307_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i307_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i307_2_NO_SHIFT_REG = rnode_168to169_bb2_add_i307_0_reg_169_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_add_i771_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i771_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i771_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i771_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i771_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i771_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_add_i771_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_add_i771_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_add_i771_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_add_i771_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_add_i771_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_add_i771_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_add_i771_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_add_i771_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_add_i771_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_168to169_bb2_add_i771_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_add_i771_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_add_i771_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_add_i771_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i771_0_stall_in_0_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i771_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i771_0_NO_SHIFT_REG = rnode_168to169_bb2_add_i771_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i771_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i771_1_NO_SHIFT_REG = rnode_168to169_bb2_add_i771_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i771_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i771_2_NO_SHIFT_REG = rnode_168to169_bb2_add_i771_0_reg_169_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_add_i399_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i399_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i399_1_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i399_2_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_168to169_bb2_add_i399_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_valid_out_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_stall_in_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_add_i399_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_add_i399_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_add_i399_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_add_i399_0_stall_in_0_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_add_i399_0_valid_out_0_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_add_i399_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_add_i399_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_add_i399_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_add_i399_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_add_i399_0_reg_169_fifo.DATA_WIDTH = 32;
defparam rnode_168to169_bb2_add_i399_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_add_i399_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_add_i399_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_add_i399_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i399_0_stall_in_0_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i399_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i399_0_NO_SHIFT_REG = rnode_168to169_bb2_add_i399_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i399_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i399_1_NO_SHIFT_REG = rnode_168to169_bb2_add_i399_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_add_i399_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_168to169_bb2_add_i399_2_NO_SHIFT_REG = rnode_168to169_bb2_add_i399_0_reg_169_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i16_i_stall_local;
wire [31:0] local_bb2_shr_i16_i;

assign local_bb2_shr_i16_i = (local_bb2_conv3_i_i >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i18_i_stall_local;
wire [31:0] local_bb2_shl1_i18_i;

assign local_bb2_shl1_i18_i = (local_bb2_conv3_i_i << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u70_stall_local;
wire [31:0] local_bb2_var__u70;

assign local_bb2_var__u70 = (local_bb2_conv3_i_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i_i_stall_local;
wire [31:0] local_bb2_shl1_i_i;

assign local_bb2_shl1_i_i = (local_bb2_conv3_i_i << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb2__tr_i_stall_local;
wire [31:0] local_bb2__tr_i;

assign local_bb2__tr_i = local_bb2_var__u62[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i16_i1408_stall_local;
wire [31:0] local_bb2_shr_i16_i1408;

assign local_bb2_shr_i16_i1408 = (local_bb2_conv3_i_i1405 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i18_i1410_stall_local;
wire [31:0] local_bb2_shl1_i18_i1410;

assign local_bb2_shl1_i18_i1410 = (local_bb2_conv3_i_i1405 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u71_stall_local;
wire [31:0] local_bb2_var__u71;

assign local_bb2_var__u71 = (local_bb2_conv3_i_i1405 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i_i1418_stall_local;
wire [31:0] local_bb2_shl1_i_i1418;

assign local_bb2_shl1_i_i1418 = (local_bb2_conv3_i_i1405 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb2__tr_i1406_stall_local;
wire [31:0] local_bb2__tr_i1406;

assign local_bb2__tr_i1406 = local_bb2_var__u63[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i16_i860_stall_local;
wire [31:0] local_bb2_shr_i16_i860;

assign local_bb2_shr_i16_i860 = (local_bb2_conv3_i_i857 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i18_i862_stall_local;
wire [31:0] local_bb2_shl1_i18_i862;

assign local_bb2_shl1_i18_i862 = (local_bb2_conv3_i_i857 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u72_stall_local;
wire [31:0] local_bb2_var__u72;

assign local_bb2_var__u72 = (local_bb2_conv3_i_i857 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i_i870_stall_local;
wire [31:0] local_bb2_shl1_i_i870;

assign local_bb2_shl1_i_i870 = (local_bb2_conv3_i_i857 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb2__tr_i858_stall_local;
wire [31:0] local_bb2__tr_i858;

assign local_bb2__tr_i858 = local_bb2_var__u64[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i16_i396_stall_local;
wire [31:0] local_bb2_shr_i16_i396;

assign local_bb2_shr_i16_i396 = (local_bb2_conv3_i_i393 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i18_i398_stall_local;
wire [31:0] local_bb2_shl1_i18_i398;

assign local_bb2_shl1_i18_i398 = (local_bb2_conv3_i_i393 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u73_stall_local;
wire [31:0] local_bb2_var__u73;

assign local_bb2_var__u73 = (local_bb2_conv3_i_i393 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i_i406_stall_local;
wire [31:0] local_bb2_shl1_i_i406;

assign local_bb2_shl1_i_i406 = (local_bb2_conv3_i_i393 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb2__tr_i394_stall_local;
wire [31:0] local_bb2__tr_i394;

assign local_bb2__tr_i394 = local_bb2_var__u65[31:0];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_reduction_0_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_reduction_0_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_reduction_0_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_reduction_0_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_reduction_0_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_reduction_0_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_reduction_0_i_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_reduction_0_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_reduction_0_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_reduction_0_i_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_reduction_0_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_reduction_0_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_reduction_0_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_reduction_0_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i_0_NO_SHIFT_REG = rnode_169to170_bb2_reduction_0_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_reduction_0_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_var__u46_0_valid_out_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u46_0_stall_in_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u46_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u46_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u46_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u46_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u46_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u46_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_var__u46_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_var__u46_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_var__u46_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_var__u46_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_var__u46_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_var__u46_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_var__u46_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_var__u46_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_var__u46_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_168to169_bb2_var__u46_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_var__u46_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_var__u46_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_var__u46_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u46_0_NO_SHIFT_REG = rnode_168to169_bb2_var__u46_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_var__u46_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u46_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_reduction_0_i1337_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1337_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1337_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1337_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1337_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1337_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1337_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1337_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_reduction_0_i1337_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_reduction_0_i1337_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_reduction_0_i1337_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_reduction_0_i1337_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_reduction_0_i1337_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_reduction_0_i1337_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_reduction_0_i1337_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_reduction_0_i1337_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_reduction_0_i1337_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_reduction_0_i1337_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_reduction_0_i1337_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_reduction_0_i1337_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_reduction_0_i1337_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1337_0_NO_SHIFT_REG = rnode_169to170_bb2_reduction_0_i1337_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_reduction_0_i1337_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1337_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_var__u56_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u56_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u56_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u56_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u56_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u56_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u56_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u56_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_var__u56_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_var__u56_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_var__u56_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_var__u56_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_var__u56_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_var__u56_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_var__u56_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_var__u56_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_var__u56_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_var__u56_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_var__u56_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_var__u56_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_var__u56_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u56_0_NO_SHIFT_REG = rnode_169to170_bb2_var__u56_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_var__u56_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u56_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i16_i1865_stall_local;
wire [31:0] local_bb2_shr_i16_i1865;

assign local_bb2_shr_i16_i1865 = (local_bb2_conv3_i_i1862 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i18_i1867_stall_local;
wire [31:0] local_bb2_shl1_i18_i1867;

assign local_bb2_shl1_i18_i1867 = (local_bb2_conv3_i_i1862 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u74_stall_local;
wire [31:0] local_bb2_var__u74;

assign local_bb2_var__u74 = (local_bb2_conv3_i_i1862 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i_i1875_stall_local;
wire [31:0] local_bb2_shl1_i_i1875;

assign local_bb2_shl1_i_i1875 = (local_bb2_conv3_i_i1862 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb2__tr_i1863_stall_local;
wire [31:0] local_bb2__tr_i1863;

assign local_bb2__tr_i1863 = local_bb2_var__u66[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i16_i1316_stall_local;
wire [31:0] local_bb2_shr_i16_i1316;

assign local_bb2_shr_i16_i1316 = (local_bb2_conv3_i_i1313 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i18_i1318_stall_local;
wire [31:0] local_bb2_shl1_i18_i1318;

assign local_bb2_shl1_i18_i1318 = (local_bb2_conv3_i_i1313 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u75_stall_local;
wire [31:0] local_bb2_var__u75;

assign local_bb2_var__u75 = (local_bb2_conv3_i_i1313 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i_i1326_stall_local;
wire [31:0] local_bb2_shl1_i_i1326;

assign local_bb2_shl1_i_i1326 = (local_bb2_conv3_i_i1313 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb2__tr_i1314_stall_local;
wire [31:0] local_bb2__tr_i1314;

assign local_bb2__tr_i1314 = local_bb2_var__u67[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i16_i768_stall_local;
wire [31:0] local_bb2_shr_i16_i768;

assign local_bb2_shr_i16_i768 = (local_bb2_conv3_i_i765 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i18_i770_stall_local;
wire [31:0] local_bb2_shl1_i18_i770;

assign local_bb2_shl1_i18_i770 = (local_bb2_conv3_i_i765 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u76_stall_local;
wire [31:0] local_bb2_var__u76;

assign local_bb2_var__u76 = (local_bb2_conv3_i_i765 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i_i778_stall_local;
wire [31:0] local_bb2_shl1_i_i778;

assign local_bb2_shl1_i_i778 = (local_bb2_conv3_i_i765 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb2__tr_i766_stall_local;
wire [31:0] local_bb2__tr_i766;

assign local_bb2__tr_i766 = local_bb2_var__u68[31:0];

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i16_i304_stall_local;
wire [31:0] local_bb2_shr_i16_i304;

assign local_bb2_shr_i16_i304 = (local_bb2_conv3_i_i301 >> 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i18_i306_stall_local;
wire [31:0] local_bb2_shl1_i18_i306;

assign local_bb2_shl1_i18_i306 = (local_bb2_conv3_i_i301 << 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u77_stall_local;
wire [31:0] local_bb2_var__u77;

assign local_bb2_var__u77 = (local_bb2_conv3_i_i301 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shl1_i_i314_stall_local;
wire [31:0] local_bb2_shl1_i_i314;

assign local_bb2_shl1_i_i314 = (local_bb2_conv3_i_i301 << 32'h9);

// This section implements an unregistered operation.
// 
wire local_bb2__tr_i302_stall_local;
wire [31:0] local_bb2__tr_i302;

assign local_bb2__tr_i302 = local_bb2_var__u69[31:0];

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_reduction_0_i1886_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1886_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1886_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1886_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1886_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1886_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1886_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1886_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_reduction_0_i1886_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_reduction_0_i1886_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_reduction_0_i1886_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_reduction_0_i1886_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_reduction_0_i1886_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_reduction_0_i1886_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_reduction_0_i1886_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_reduction_0_i1886_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_reduction_0_i1886_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_reduction_0_i1886_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_reduction_0_i1886_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_reduction_0_i1886_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_reduction_0_i1886_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1886_0_NO_SHIFT_REG = rnode_169to170_bb2_reduction_0_i1886_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_reduction_0_i1886_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1886_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_var__u54_0_valid_out_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u54_0_stall_in_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u54_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u54_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u54_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u54_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u54_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u54_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_var__u54_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_var__u54_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_var__u54_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_var__u54_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_var__u54_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_var__u54_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_var__u54_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_var__u54_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_var__u54_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_168to169_bb2_var__u54_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_var__u54_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_var__u54_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_var__u54_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u54_0_NO_SHIFT_REG = rnode_168to169_bb2_var__u54_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_var__u54_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u54_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_reduction_0_i1429_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1429_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1429_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1429_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1429_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1429_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1429_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i1429_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_reduction_0_i1429_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_reduction_0_i1429_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_reduction_0_i1429_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_reduction_0_i1429_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_reduction_0_i1429_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_reduction_0_i1429_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_reduction_0_i1429_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_reduction_0_i1429_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_reduction_0_i1429_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_reduction_0_i1429_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_reduction_0_i1429_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_reduction_0_i1429_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_reduction_0_i1429_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1429_0_NO_SHIFT_REG = rnode_169to170_bb2_reduction_0_i1429_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_reduction_0_i1429_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1429_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_var__u48_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u48_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u48_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u48_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u48_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u48_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u48_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u48_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_var__u48_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_var__u48_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_var__u48_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_var__u48_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_var__u48_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_var__u48_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_var__u48_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_var__u48_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_var__u48_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_var__u48_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_var__u48_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_var__u48_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_var__u48_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u48_0_NO_SHIFT_REG = rnode_169to170_bb2_var__u48_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_var__u48_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u48_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_reduction_0_i881_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i881_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i881_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i881_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i881_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i881_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i881_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i881_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_reduction_0_i881_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_reduction_0_i881_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_reduction_0_i881_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_reduction_0_i881_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_reduction_0_i881_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_reduction_0_i881_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_reduction_0_i881_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_reduction_0_i881_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_reduction_0_i881_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_reduction_0_i881_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_reduction_0_i881_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_reduction_0_i881_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_reduction_0_i881_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i881_0_NO_SHIFT_REG = rnode_169to170_bb2_reduction_0_i881_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_reduction_0_i881_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i881_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_var__u50_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u50_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u50_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u50_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u50_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u50_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u50_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u50_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_var__u50_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_var__u50_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_var__u50_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_var__u50_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_var__u50_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_var__u50_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_var__u50_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_var__u50_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_var__u50_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_var__u50_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_var__u50_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_var__u50_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_var__u50_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u50_0_NO_SHIFT_REG = rnode_169to170_bb2_var__u50_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_var__u50_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u50_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_reduction_0_i325_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i325_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i325_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i325_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i325_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i325_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i325_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i325_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_reduction_0_i325_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_reduction_0_i325_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_reduction_0_i325_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_reduction_0_i325_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_reduction_0_i325_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_reduction_0_i325_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_reduction_0_i325_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_reduction_0_i325_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_reduction_0_i325_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_reduction_0_i325_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_reduction_0_i325_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_reduction_0_i325_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_reduction_0_i325_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i325_0_NO_SHIFT_REG = rnode_169to170_bb2_reduction_0_i325_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_reduction_0_i325_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i325_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_var__u60_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u60_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u60_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u60_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u60_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u60_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u60_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u60_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_var__u60_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_var__u60_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_var__u60_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_var__u60_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_var__u60_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_var__u60_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_var__u60_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_var__u60_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_var__u60_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_var__u60_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_var__u60_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_var__u60_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_var__u60_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u60_0_NO_SHIFT_REG = rnode_169to170_bb2_var__u60_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_var__u60_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u60_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_reduction_0_i789_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i789_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i789_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i789_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i789_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i789_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i789_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i789_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_reduction_0_i789_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_reduction_0_i789_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_reduction_0_i789_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_reduction_0_i789_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_reduction_0_i789_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_reduction_0_i789_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_reduction_0_i789_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_reduction_0_i789_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_reduction_0_i789_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_reduction_0_i789_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_reduction_0_i789_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_reduction_0_i789_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_reduction_0_i789_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i789_0_NO_SHIFT_REG = rnode_169to170_bb2_reduction_0_i789_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_reduction_0_i789_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i789_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_168to169_bb2_var__u58_0_valid_out_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u58_0_stall_in_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u58_0_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u58_0_reg_169_inputs_ready_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u58_0_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u58_0_valid_out_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u58_0_stall_in_reg_169_NO_SHIFT_REG;
 logic rnode_168to169_bb2_var__u58_0_stall_out_reg_169_NO_SHIFT_REG;

acl_data_fifo rnode_168to169_bb2_var__u58_0_reg_169_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_168to169_bb2_var__u58_0_reg_169_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_168to169_bb2_var__u58_0_stall_in_reg_169_NO_SHIFT_REG),
	.valid_out(rnode_168to169_bb2_var__u58_0_valid_out_reg_169_NO_SHIFT_REG),
	.stall_out(rnode_168to169_bb2_var__u58_0_stall_out_reg_169_NO_SHIFT_REG),
	.data_in(rnode_167to168_bb2_var__u58_0_NO_SHIFT_REG),
	.data_out(rnode_168to169_bb2_var__u58_0_reg_169_NO_SHIFT_REG)
);

defparam rnode_168to169_bb2_var__u58_0_reg_169_fifo.DEPTH = 1;
defparam rnode_168to169_bb2_var__u58_0_reg_169_fifo.DATA_WIDTH = 1;
defparam rnode_168to169_bb2_var__u58_0_reg_169_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_168to169_bb2_var__u58_0_reg_169_fifo.IMPL = "shift_reg";

assign rnode_168to169_bb2_var__u58_0_reg_169_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to168_bb2_var__u58_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u58_0_NO_SHIFT_REG = rnode_168to169_bb2_var__u58_0_reg_169_NO_SHIFT_REG;
assign rnode_168to169_bb2_var__u58_0_stall_in_reg_169_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u58_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_reduction_0_i417_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i417_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i417_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i417_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i417_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i417_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i417_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_reduction_0_i417_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_reduction_0_i417_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_reduction_0_i417_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_reduction_0_i417_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_reduction_0_i417_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_reduction_0_i417_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_reduction_0_i417_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_reduction_0_i417_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_reduction_0_i417_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_reduction_0_i417_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_reduction_0_i417_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_reduction_0_i417_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_reduction_0_i417_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_reduction_0_i417_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i417_0_NO_SHIFT_REG = rnode_169to170_bb2_reduction_0_i417_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_reduction_0_i417_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i417_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_var__u52_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u52_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u52_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u52_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u52_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u52_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u52_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_var__u52_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_var__u52_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_var__u52_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_var__u52_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_var__u52_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_var__u52_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2_var__u52_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2_var__u52_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_var__u52_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_var__u52_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_var__u52_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_var__u52_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_var__u52_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2_var__u52_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u52_0_NO_SHIFT_REG = rnode_169to170_bb2_var__u52_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_var__u52_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u52_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__29_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__29_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__29_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__29_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__29_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__29_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2__29_i_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2__29_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__29_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__29_i_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__29_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__29_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__29_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2__29_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i_0_NO_SHIFT_REG = rnode_169to170_bb2__29_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__29_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__29_i1399_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1399_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1399_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1399_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1399_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1399_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1399_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1399_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__29_i1399_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__29_i1399_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__29_i1399_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__29_i1399_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__29_i1399_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2__29_i1399_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2__29_i1399_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__29_i1399_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__29_i1399_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__29_i1399_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__29_i1399_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__29_i1399_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2__29_i1399_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1399_0_NO_SHIFT_REG = rnode_169to170_bb2__29_i1399_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__29_i1399_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1399_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__29_i851_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i851_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i851_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i851_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i851_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i851_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i851_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i851_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__29_i851_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__29_i851_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__29_i851_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__29_i851_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__29_i851_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2__29_i851_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2__29_i851_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__29_i851_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__29_i851_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__29_i851_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__29_i851_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__29_i851_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2__29_i851_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i851_0_NO_SHIFT_REG = rnode_169to170_bb2__29_i851_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__29_i851_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i851_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__29_i387_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i387_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i387_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i387_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i387_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i387_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i387_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i387_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__29_i387_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__29_i387_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__29_i387_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__29_i387_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__29_i387_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2__29_i387_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2__29_i387_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__29_i387_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__29_i387_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__29_i387_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__29_i387_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__29_i387_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2__29_i387_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i387_0_NO_SHIFT_REG = rnode_169to170_bb2__29_i387_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__29_i387_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i387_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__29_i1307_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1307_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1307_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1307_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1307_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1307_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1307_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1307_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__29_i1307_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__29_i1307_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__29_i1307_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__29_i1307_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__29_i1307_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2__29_i1307_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2__29_i1307_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__29_i1307_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__29_i1307_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__29_i1307_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__29_i1307_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__29_i1307_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2__29_i1307_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1307_0_NO_SHIFT_REG = rnode_169to170_bb2__29_i1307_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__29_i1307_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1307_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__29_i1856_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1856_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1856_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1856_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1856_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1856_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1856_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i1856_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__29_i1856_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__29_i1856_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__29_i1856_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__29_i1856_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__29_i1856_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2__29_i1856_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2__29_i1856_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__29_i1856_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__29_i1856_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__29_i1856_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__29_i1856_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__29_i1856_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2__29_i1856_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1856_0_NO_SHIFT_REG = rnode_169to170_bb2__29_i1856_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__29_i1856_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1856_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__29_i759_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i759_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i759_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i759_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i759_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i759_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i759_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i759_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__29_i759_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__29_i759_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__29_i759_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__29_i759_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__29_i759_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2__29_i759_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2__29_i759_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__29_i759_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__29_i759_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__29_i759_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__29_i759_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__29_i759_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2__29_i759_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i759_0_NO_SHIFT_REG = rnode_169to170_bb2__29_i759_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__29_i759_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i759_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__29_i295_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i295_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i295_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i295_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i295_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i295_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i295_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__29_i295_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__29_i295_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__29_i295_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__29_i295_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__29_i295_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__29_i295_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(rnode_167to169_bb2__29_i295_0_NO_SHIFT_REG),
	.data_out(rnode_169to170_bb2__29_i295_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__29_i295_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__29_i295_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__29_i295_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__29_i295_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__29_i295_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_167to169_bb2__29_i295_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i295_0_NO_SHIFT_REG = rnode_169to170_bb2__29_i295_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__29_i295_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i295_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and4_i_stall_local;
wire [31:0] local_bb2_and4_i;

assign local_bb2_and4_i = (rnode_169to170_bb2_xor_i_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and4_i1279_stall_local;
wire [31:0] local_bb2_and4_i1279;

assign local_bb2_and4_i1279 = (rnode_169to170_bb2_xor_i1278_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and4_i1828_stall_local;
wire [31:0] local_bb2_and4_i1828;

assign local_bb2_and4_i1828 = (rnode_169to170_bb2_xor_i1827_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and4_i1371_stall_local;
wire [31:0] local_bb2_and4_i1371;

assign local_bb2_and4_i1371 = (rnode_169to170_bb2_xor_i1370_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and4_i823_stall_local;
wire [31:0] local_bb2_and4_i823;

assign local_bb2_and4_i823 = (rnode_169to170_bb2_xor_i822_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and4_i267_stall_local;
wire [31:0] local_bb2_and4_i267;

assign local_bb2_and4_i267 = (rnode_169to170_bb2_xor_i266_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and4_i731_stall_local;
wire [31:0] local_bb2_and4_i731;

assign local_bb2_and4_i731 = (rnode_169to170_bb2_xor_i730_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and4_i359_stall_local;
wire [31:0] local_bb2_and4_i359;

assign local_bb2_and4_i359 = (rnode_169to170_bb2_xor_i358_0_NO_SHIFT_REG & 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_inc_i_stall_local;
wire [31:0] local_bb2_inc_i;

assign local_bb2_inc_i = (rnode_168to169_bb2_add_i_0_NO_SHIFT_REG + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp50_not_i_stall_local;
wire local_bb2_cmp50_not_i;

assign local_bb2_cmp50_not_i = (rnode_168to169_bb2_add_i_1_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_inc_i1322_stall_local;
wire [31:0] local_bb2_inc_i1322;

assign local_bb2_inc_i1322 = (rnode_168to169_bb2_add_i1319_0_NO_SHIFT_REG + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp50_not_i1327_stall_local;
wire local_bb2_cmp50_not_i1327;

assign local_bb2_cmp50_not_i1327 = (rnode_168to169_bb2_add_i1319_1_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_inc_i1871_stall_local;
wire [31:0] local_bb2_inc_i1871;

assign local_bb2_inc_i1871 = (rnode_168to169_bb2_add_i1868_0_NO_SHIFT_REG + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp50_not_i1876_stall_local;
wire local_bb2_cmp50_not_i1876;

assign local_bb2_cmp50_not_i1876 = (rnode_168to169_bb2_add_i1868_1_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_inc_i1414_stall_local;
wire [31:0] local_bb2_inc_i1414;

assign local_bb2_inc_i1414 = (rnode_168to169_bb2_add_i1411_0_NO_SHIFT_REG + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp50_not_i1419_stall_local;
wire local_bb2_cmp50_not_i1419;

assign local_bb2_cmp50_not_i1419 = (rnode_168to169_bb2_add_i1411_1_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_inc_i866_stall_local;
wire [31:0] local_bb2_inc_i866;

assign local_bb2_inc_i866 = (rnode_168to169_bb2_add_i863_0_NO_SHIFT_REG + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp50_not_i871_stall_local;
wire local_bb2_cmp50_not_i871;

assign local_bb2_cmp50_not_i871 = (rnode_168to169_bb2_add_i863_1_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_inc_i310_stall_local;
wire [31:0] local_bb2_inc_i310;

assign local_bb2_inc_i310 = (rnode_168to169_bb2_add_i307_0_NO_SHIFT_REG + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp50_not_i315_stall_local;
wire local_bb2_cmp50_not_i315;

assign local_bb2_cmp50_not_i315 = (rnode_168to169_bb2_add_i307_1_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_inc_i774_stall_local;
wire [31:0] local_bb2_inc_i774;

assign local_bb2_inc_i774 = (rnode_168to169_bb2_add_i771_0_NO_SHIFT_REG + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp50_not_i779_stall_local;
wire local_bb2_cmp50_not_i779;

assign local_bb2_cmp50_not_i779 = (rnode_168to169_bb2_add_i771_1_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_inc_i402_stall_local;
wire [31:0] local_bb2_inc_i402;

assign local_bb2_inc_i402 = (rnode_168to169_bb2_add_i399_0_NO_SHIFT_REG + 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp50_not_i407_stall_local;
wire local_bb2_cmp50_not_i407;

assign local_bb2_cmp50_not_i407 = (rnode_168to169_bb2_add_i399_1_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i_stall_local;
wire [31:0] local_bb2_shr_i_i;

assign local_bb2_shr_i_i = (local_bb2_var__u70 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i15_i_stall_local;
wire [31:0] local_bb2_shl_i15_i;

assign local_bb2_shl_i15_i = (local_bb2__tr_i & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and48_i_stall_local;
wire [31:0] local_bb2_and48_i;

assign local_bb2_and48_i = (local_bb2__tr_i & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i1416_stall_local;
wire [31:0] local_bb2_shr_i_i1416;

assign local_bb2_shr_i_i1416 = (local_bb2_var__u71 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i15_i1407_stall_local;
wire [31:0] local_bb2_shl_i15_i1407;

assign local_bb2_shl_i15_i1407 = (local_bb2__tr_i1406 & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and48_i1412_stall_local;
wire [31:0] local_bb2_and48_i1412;

assign local_bb2_and48_i1412 = (local_bb2__tr_i1406 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i868_stall_local;
wire [31:0] local_bb2_shr_i_i868;

assign local_bb2_shr_i_i868 = (local_bb2_var__u72 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i15_i859_stall_local;
wire [31:0] local_bb2_shl_i15_i859;

assign local_bb2_shl_i15_i859 = (local_bb2__tr_i858 & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and48_i864_stall_local;
wire [31:0] local_bb2_and48_i864;

assign local_bb2_and48_i864 = (local_bb2__tr_i858 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i404_stall_local;
wire [31:0] local_bb2_shr_i_i404;

assign local_bb2_shr_i_i404 = (local_bb2_var__u73 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i15_i395_stall_local;
wire [31:0] local_bb2_shl_i15_i395;

assign local_bb2_shl_i15_i395 = (local_bb2__tr_i394 & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and48_i400_stall_local;
wire [31:0] local_bb2_and48_i400;

assign local_bb2_and48_i400 = (local_bb2__tr_i394 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i1873_stall_local;
wire [31:0] local_bb2_shr_i_i1873;

assign local_bb2_shr_i_i1873 = (local_bb2_var__u74 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i15_i1864_stall_local;
wire [31:0] local_bb2_shl_i15_i1864;

assign local_bb2_shl_i15_i1864 = (local_bb2__tr_i1863 & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and48_i1869_stall_local;
wire [31:0] local_bb2_and48_i1869;

assign local_bb2_and48_i1869 = (local_bb2__tr_i1863 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i1324_stall_local;
wire [31:0] local_bb2_shr_i_i1324;

assign local_bb2_shr_i_i1324 = (local_bb2_var__u75 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i15_i1315_stall_local;
wire [31:0] local_bb2_shl_i15_i1315;

assign local_bb2_shl_i15_i1315 = (local_bb2__tr_i1314 & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and48_i1320_stall_local;
wire [31:0] local_bb2_and48_i1320;

assign local_bb2_and48_i1320 = (local_bb2__tr_i1314 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i776_stall_local;
wire [31:0] local_bb2_shr_i_i776;

assign local_bb2_shr_i_i776 = (local_bb2_var__u76 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i15_i767_stall_local;
wire [31:0] local_bb2_shl_i15_i767;

assign local_bb2_shl_i15_i767 = (local_bb2__tr_i766 & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and48_i772_stall_local;
wire [31:0] local_bb2_and48_i772;

assign local_bb2_and48_i772 = (local_bb2__tr_i766 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i312_stall_local;
wire [31:0] local_bb2_shr_i_i312;

assign local_bb2_shr_i_i312 = (local_bb2_var__u77 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i15_i303_stall_local;
wire [31:0] local_bb2_shl_i15_i303;

assign local_bb2_shl_i15_i303 = (local_bb2__tr_i302 & 32'hFFFF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and48_i308_stall_local;
wire [31:0] local_bb2_and48_i308;

assign local_bb2_and48_i308 = (local_bb2__tr_i302 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i17_i_stall_local;
wire [31:0] local_bb2_or_i17_i;

assign local_bb2_or_i17_i = (local_bb2_shl_i15_i | local_bb2_shr_i16_i);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool49_i_stall_local;
wire local_bb2_tobool49_i;

assign local_bb2_tobool49_i = (local_bb2_and48_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i17_i1409_stall_local;
wire [31:0] local_bb2_or_i17_i1409;

assign local_bb2_or_i17_i1409 = (local_bb2_shl_i15_i1407 | local_bb2_shr_i16_i1408);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool49_i1413_stall_local;
wire local_bb2_tobool49_i1413;

assign local_bb2_tobool49_i1413 = (local_bb2_and48_i1412 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i17_i861_stall_local;
wire [31:0] local_bb2_or_i17_i861;

assign local_bb2_or_i17_i861 = (local_bb2_shl_i15_i859 | local_bb2_shr_i16_i860);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool49_i865_stall_local;
wire local_bb2_tobool49_i865;

assign local_bb2_tobool49_i865 = (local_bb2_and48_i864 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i17_i397_stall_local;
wire [31:0] local_bb2_or_i17_i397;

assign local_bb2_or_i17_i397 = (local_bb2_shl_i15_i395 | local_bb2_shr_i16_i396);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool49_i401_stall_local;
wire local_bb2_tobool49_i401;

assign local_bb2_tobool49_i401 = (local_bb2_and48_i400 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i17_i1866_stall_local;
wire [31:0] local_bb2_or_i17_i1866;

assign local_bb2_or_i17_i1866 = (local_bb2_shl_i15_i1864 | local_bb2_shr_i16_i1865);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool49_i1870_stall_local;
wire local_bb2_tobool49_i1870;

assign local_bb2_tobool49_i1870 = (local_bb2_and48_i1869 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i17_i1317_stall_local;
wire [31:0] local_bb2_or_i17_i1317;

assign local_bb2_or_i17_i1317 = (local_bb2_shl_i15_i1315 | local_bb2_shr_i16_i1316);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool49_i1321_stall_local;
wire local_bb2_tobool49_i1321;

assign local_bb2_tobool49_i1321 = (local_bb2_and48_i1320 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i17_i769_stall_local;
wire [31:0] local_bb2_or_i17_i769;

assign local_bb2_or_i17_i769 = (local_bb2_shl_i15_i767 | local_bb2_shr_i16_i768);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool49_i773_stall_local;
wire local_bb2_tobool49_i773;

assign local_bb2_tobool49_i773 = (local_bb2_and48_i772 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i17_i305_stall_local;
wire [31:0] local_bb2_or_i17_i305;

assign local_bb2_or_i17_i305 = (local_bb2_shl_i15_i303 | local_bb2_shr_i16_i304);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool49_i309_stall_local;
wire local_bb2_tobool49_i309;

assign local_bb2_tobool49_i309 = (local_bb2_and48_i308 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_i_stall_local;
wire [31:0] local_bb2_shl_i_i;

assign local_bb2_shl_i_i = (local_bb2_or_i17_i << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i_stall_local;
wire local_bb2__31_i;

assign local_bb2__31_i = (local_bb2_tobool49_i & local_bb2_cmp50_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_i1415_stall_local;
wire [31:0] local_bb2_shl_i_i1415;

assign local_bb2_shl_i_i1415 = (local_bb2_or_i17_i1409 << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i1420_stall_local;
wire local_bb2__31_i1420;

assign local_bb2__31_i1420 = (local_bb2_tobool49_i1413 & local_bb2_cmp50_not_i1419);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_i867_stall_local;
wire [31:0] local_bb2_shl_i_i867;

assign local_bb2_shl_i_i867 = (local_bb2_or_i17_i861 << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i872_stall_local;
wire local_bb2__31_i872;

assign local_bb2__31_i872 = (local_bb2_tobool49_i865 & local_bb2_cmp50_not_i871);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_i403_stall_local;
wire [31:0] local_bb2_shl_i_i403;

assign local_bb2_shl_i_i403 = (local_bb2_or_i17_i397 << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i408_stall_local;
wire local_bb2__31_i408;

assign local_bb2__31_i408 = (local_bb2_tobool49_i401 & local_bb2_cmp50_not_i407);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_i1872_stall_local;
wire [31:0] local_bb2_shl_i_i1872;

assign local_bb2_shl_i_i1872 = (local_bb2_or_i17_i1866 << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i1877_stall_local;
wire local_bb2__31_i1877;

assign local_bb2__31_i1877 = (local_bb2_tobool49_i1870 & local_bb2_cmp50_not_i1876);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_i1323_stall_local;
wire [31:0] local_bb2_shl_i_i1323;

assign local_bb2_shl_i_i1323 = (local_bb2_or_i17_i1317 << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i1328_stall_local;
wire local_bb2__31_i1328;

assign local_bb2__31_i1328 = (local_bb2_tobool49_i1321 & local_bb2_cmp50_not_i1327);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_i775_stall_local;
wire [31:0] local_bb2_shl_i_i775;

assign local_bb2_shl_i_i775 = (local_bb2_or_i17_i769 << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i780_stall_local;
wire local_bb2__31_i780;

assign local_bb2__31_i780 = (local_bb2_tobool49_i773 & local_bb2_cmp50_not_i779);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_i311_stall_local;
wire [31:0] local_bb2_shl_i_i311;

assign local_bb2_shl_i_i311 = (local_bb2_or_i17_i305 << 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i316_stall_local;
wire local_bb2__31_i316;

assign local_bb2__31_i316 = (local_bb2_tobool49_i309 & local_bb2_cmp50_not_i315);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i_stall_local;
wire [31:0] local_bb2_or_i_i;

assign local_bb2_or_i_i = (local_bb2_shl_i_i | local_bb2_shr_i_i);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i_stall_local;
wire [31:0] local_bb2__32_i;

assign local_bb2__32_i = (local_bb2__31_i ? local_bb2_shl1_i_i : local_bb2_shl1_i18_i);

// This section implements an unregistered operation.
// 
wire local_bb2__36_i_stall_local;
wire [31:0] local_bb2__36_i;

assign local_bb2__36_i = (local_bb2__31_i ? rnode_168to169_bb2_add_i_2_NO_SHIFT_REG : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i1417_stall_local;
wire [31:0] local_bb2_or_i_i1417;

assign local_bb2_or_i_i1417 = (local_bb2_shl_i_i1415 | local_bb2_shr_i_i1416);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i1421_stall_local;
wire [31:0] local_bb2__32_i1421;

assign local_bb2__32_i1421 = (local_bb2__31_i1420 ? local_bb2_shl1_i_i1418 : local_bb2_shl1_i18_i1410);

// This section implements an unregistered operation.
// 
wire local_bb2__36_i1425_stall_local;
wire [31:0] local_bb2__36_i1425;

assign local_bb2__36_i1425 = (local_bb2__31_i1420 ? rnode_168to169_bb2_add_i1411_2_NO_SHIFT_REG : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i869_stall_local;
wire [31:0] local_bb2_or_i_i869;

assign local_bb2_or_i_i869 = (local_bb2_shl_i_i867 | local_bb2_shr_i_i868);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i873_stall_local;
wire [31:0] local_bb2__32_i873;

assign local_bb2__32_i873 = (local_bb2__31_i872 ? local_bb2_shl1_i_i870 : local_bb2_shl1_i18_i862);

// This section implements an unregistered operation.
// 
wire local_bb2__36_i877_stall_local;
wire [31:0] local_bb2__36_i877;

assign local_bb2__36_i877 = (local_bb2__31_i872 ? rnode_168to169_bb2_add_i863_2_NO_SHIFT_REG : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i405_stall_local;
wire [31:0] local_bb2_or_i_i405;

assign local_bb2_or_i_i405 = (local_bb2_shl_i_i403 | local_bb2_shr_i_i404);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i409_stall_local;
wire [31:0] local_bb2__32_i409;

assign local_bb2__32_i409 = (local_bb2__31_i408 ? local_bb2_shl1_i_i406 : local_bb2_shl1_i18_i398);

// This section implements an unregistered operation.
// 
wire local_bb2__36_i413_stall_local;
wire [31:0] local_bb2__36_i413;

assign local_bb2__36_i413 = (local_bb2__31_i408 ? rnode_168to169_bb2_add_i399_2_NO_SHIFT_REG : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i1874_stall_local;
wire [31:0] local_bb2_or_i_i1874;

assign local_bb2_or_i_i1874 = (local_bb2_shl_i_i1872 | local_bb2_shr_i_i1873);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i1878_stall_local;
wire [31:0] local_bb2__32_i1878;

assign local_bb2__32_i1878 = (local_bb2__31_i1877 ? local_bb2_shl1_i_i1875 : local_bb2_shl1_i18_i1867);

// This section implements an unregistered operation.
// 
wire local_bb2__36_i1882_stall_local;
wire [31:0] local_bb2__36_i1882;

assign local_bb2__36_i1882 = (local_bb2__31_i1877 ? rnode_168to169_bb2_add_i1868_2_NO_SHIFT_REG : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i1325_stall_local;
wire [31:0] local_bb2_or_i_i1325;

assign local_bb2_or_i_i1325 = (local_bb2_shl_i_i1323 | local_bb2_shr_i_i1324);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i1329_stall_local;
wire [31:0] local_bb2__32_i1329;

assign local_bb2__32_i1329 = (local_bb2__31_i1328 ? local_bb2_shl1_i_i1326 : local_bb2_shl1_i18_i1318);

// This section implements an unregistered operation.
// 
wire local_bb2__36_i1333_stall_local;
wire [31:0] local_bb2__36_i1333;

assign local_bb2__36_i1333 = (local_bb2__31_i1328 ? rnode_168to169_bb2_add_i1319_2_NO_SHIFT_REG : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i777_stall_local;
wire [31:0] local_bb2_or_i_i777;

assign local_bb2_or_i_i777 = (local_bb2_shl_i_i775 | local_bb2_shr_i_i776);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i781_stall_local;
wire [31:0] local_bb2__32_i781;

assign local_bb2__32_i781 = (local_bb2__31_i780 ? local_bb2_shl1_i_i778 : local_bb2_shl1_i18_i770);

// This section implements an unregistered operation.
// 
wire local_bb2__36_i785_stall_local;
wire [31:0] local_bb2__36_i785;

assign local_bb2__36_i785 = (local_bb2__31_i780 ? rnode_168to169_bb2_add_i771_2_NO_SHIFT_REG : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i313_stall_local;
wire [31:0] local_bb2_or_i_i313;

assign local_bb2_or_i_i313 = (local_bb2_shl_i_i311 | local_bb2_shr_i_i312);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i317_stall_local;
wire [31:0] local_bb2__32_i317;

assign local_bb2__32_i317 = (local_bb2__31_i316 ? local_bb2_shl1_i_i314 : local_bb2_shl1_i18_i306);

// This section implements an unregistered operation.
// 
wire local_bb2__36_i321_stall_local;
wire [31:0] local_bb2__36_i321;

assign local_bb2__36_i321 = (local_bb2__31_i316 ? rnode_168to169_bb2_add_i307_2_NO_SHIFT_REG : 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__34_i_stall_local;
wire [31:0] local_bb2__34_i;

assign local_bb2__34_i = (local_bb2__31_i ? local_bb2_or_i_i : local_bb2_or_i17_i);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i_stall_local;
wire [31:0] local_bb2__33_i;

assign local_bb2__33_i = (local_bb2_tobool49_i ? local_bb2__32_i : local_bb2_shl1_i18_i);

// This section implements an unregistered operation.
// 
wire local_bb2__37_i_stall_local;
wire [31:0] local_bb2__37_i;

assign local_bb2__37_i = (local_bb2_tobool49_i ? local_bb2__36_i : local_bb2_inc_i);

// This section implements an unregistered operation.
// 
wire local_bb2__34_i1423_stall_local;
wire [31:0] local_bb2__34_i1423;

assign local_bb2__34_i1423 = (local_bb2__31_i1420 ? local_bb2_or_i_i1417 : local_bb2_or_i17_i1409);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i1422_stall_local;
wire [31:0] local_bb2__33_i1422;

assign local_bb2__33_i1422 = (local_bb2_tobool49_i1413 ? local_bb2__32_i1421 : local_bb2_shl1_i18_i1410);

// This section implements an unregistered operation.
// 
wire local_bb2__37_i1426_stall_local;
wire [31:0] local_bb2__37_i1426;

assign local_bb2__37_i1426 = (local_bb2_tobool49_i1413 ? local_bb2__36_i1425 : local_bb2_inc_i1414);

// This section implements an unregistered operation.
// 
wire local_bb2__34_i875_stall_local;
wire [31:0] local_bb2__34_i875;

assign local_bb2__34_i875 = (local_bb2__31_i872 ? local_bb2_or_i_i869 : local_bb2_or_i17_i861);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i874_stall_local;
wire [31:0] local_bb2__33_i874;

assign local_bb2__33_i874 = (local_bb2_tobool49_i865 ? local_bb2__32_i873 : local_bb2_shl1_i18_i862);

// This section implements an unregistered operation.
// 
wire local_bb2__37_i878_stall_local;
wire [31:0] local_bb2__37_i878;

assign local_bb2__37_i878 = (local_bb2_tobool49_i865 ? local_bb2__36_i877 : local_bb2_inc_i866);

// This section implements an unregistered operation.
// 
wire local_bb2__34_i411_stall_local;
wire [31:0] local_bb2__34_i411;

assign local_bb2__34_i411 = (local_bb2__31_i408 ? local_bb2_or_i_i405 : local_bb2_or_i17_i397);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i410_stall_local;
wire [31:0] local_bb2__33_i410;

assign local_bb2__33_i410 = (local_bb2_tobool49_i401 ? local_bb2__32_i409 : local_bb2_shl1_i18_i398);

// This section implements an unregistered operation.
// 
wire local_bb2__37_i414_stall_local;
wire [31:0] local_bb2__37_i414;

assign local_bb2__37_i414 = (local_bb2_tobool49_i401 ? local_bb2__36_i413 : local_bb2_inc_i402);

// This section implements an unregistered operation.
// 
wire local_bb2__34_i1880_stall_local;
wire [31:0] local_bb2__34_i1880;

assign local_bb2__34_i1880 = (local_bb2__31_i1877 ? local_bb2_or_i_i1874 : local_bb2_or_i17_i1866);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i1879_stall_local;
wire [31:0] local_bb2__33_i1879;

assign local_bb2__33_i1879 = (local_bb2_tobool49_i1870 ? local_bb2__32_i1878 : local_bb2_shl1_i18_i1867);

// This section implements an unregistered operation.
// 
wire local_bb2__37_i1883_stall_local;
wire [31:0] local_bb2__37_i1883;

assign local_bb2__37_i1883 = (local_bb2_tobool49_i1870 ? local_bb2__36_i1882 : local_bb2_inc_i1871);

// This section implements an unregistered operation.
// 
wire local_bb2__34_i1331_stall_local;
wire [31:0] local_bb2__34_i1331;

assign local_bb2__34_i1331 = (local_bb2__31_i1328 ? local_bb2_or_i_i1325 : local_bb2_or_i17_i1317);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i1330_stall_local;
wire [31:0] local_bb2__33_i1330;

assign local_bb2__33_i1330 = (local_bb2_tobool49_i1321 ? local_bb2__32_i1329 : local_bb2_shl1_i18_i1318);

// This section implements an unregistered operation.
// 
wire local_bb2__37_i1334_stall_local;
wire [31:0] local_bb2__37_i1334;

assign local_bb2__37_i1334 = (local_bb2_tobool49_i1321 ? local_bb2__36_i1333 : local_bb2_inc_i1322);

// This section implements an unregistered operation.
// 
wire local_bb2__34_i783_stall_local;
wire [31:0] local_bb2__34_i783;

assign local_bb2__34_i783 = (local_bb2__31_i780 ? local_bb2_or_i_i777 : local_bb2_or_i17_i769);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i782_stall_local;
wire [31:0] local_bb2__33_i782;

assign local_bb2__33_i782 = (local_bb2_tobool49_i773 ? local_bb2__32_i781 : local_bb2_shl1_i18_i770);

// This section implements an unregistered operation.
// 
wire local_bb2__37_i786_stall_local;
wire [31:0] local_bb2__37_i786;

assign local_bb2__37_i786 = (local_bb2_tobool49_i773 ? local_bb2__36_i785 : local_bb2_inc_i774);

// This section implements an unregistered operation.
// 
wire local_bb2__34_i319_stall_local;
wire [31:0] local_bb2__34_i319;

assign local_bb2__34_i319 = (local_bb2__31_i316 ? local_bb2_or_i_i313 : local_bb2_or_i17_i305);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i318_stall_local;
wire [31:0] local_bb2__33_i318;

assign local_bb2__33_i318 = (local_bb2_tobool49_i309 ? local_bb2__32_i317 : local_bb2_shl1_i18_i306);

// This section implements an unregistered operation.
// 
wire local_bb2__37_i322_stall_local;
wire [31:0] local_bb2__37_i322;

assign local_bb2__37_i322 = (local_bb2_tobool49_i309 ? local_bb2__36_i321 : local_bb2_inc_i310);

// This section implements an unregistered operation.
// 
wire local_bb2__35_i_stall_local;
wire [31:0] local_bb2__35_i;

assign local_bb2__35_i = (local_bb2_tobool49_i ? local_bb2__34_i : local_bb2_or_i17_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i_stall_local;
wire local_bb2_cmp77_i;

assign local_bb2_cmp77_i = (local_bb2__33_i > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u78_stall_local;
wire local_bb2_var__u78;

assign local_bb2_var__u78 = ($signed(local_bb2__33_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_cmp53_i_stall_local;
wire local_bb2_cmp53_i;

assign local_bb2_cmp53_i = (local_bb2__37_i > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp68_i_stall_local;
wire local_bb2_cmp68_i;

assign local_bb2_cmp68_i = (local_bb2__37_i < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i_stall_local;
wire [31:0] local_bb2_sub_i;

assign local_bb2_sub_i = (local_bb2__37_i << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp71_not_i_stall_local;
wire local_bb2_cmp71_not_i;

assign local_bb2_cmp71_not_i = (local_bb2__37_i != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__35_i1424_stall_local;
wire [31:0] local_bb2__35_i1424;

assign local_bb2__35_i1424 = (local_bb2_tobool49_i1413 ? local_bb2__34_i1423 : local_bb2_or_i17_i1409);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i1437_stall_local;
wire local_bb2_cmp77_i1437;

assign local_bb2_cmp77_i1437 = (local_bb2__33_i1422 > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u79_stall_local;
wire local_bb2_var__u79;

assign local_bb2_var__u79 = ($signed(local_bb2__33_i1422) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2__35_i876_stall_local;
wire [31:0] local_bb2__35_i876;

assign local_bb2__35_i876 = (local_bb2_tobool49_i865 ? local_bb2__34_i875 : local_bb2_or_i17_i861);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i889_stall_local;
wire local_bb2_cmp77_i889;

assign local_bb2_cmp77_i889 = (local_bb2__33_i874 > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u80_stall_local;
wire local_bb2_var__u80;

assign local_bb2_var__u80 = ($signed(local_bb2__33_i874) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2__35_i412_stall_local;
wire [31:0] local_bb2__35_i412;

assign local_bb2__35_i412 = (local_bb2_tobool49_i401 ? local_bb2__34_i411 : local_bb2_or_i17_i397);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i425_stall_local;
wire local_bb2_cmp77_i425;

assign local_bb2_cmp77_i425 = (local_bb2__33_i410 > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u81_stall_local;
wire local_bb2_var__u81;

assign local_bb2_var__u81 = ($signed(local_bb2__33_i410) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2__35_i1881_stall_local;
wire [31:0] local_bb2__35_i1881;

assign local_bb2__35_i1881 = (local_bb2_tobool49_i1870 ? local_bb2__34_i1880 : local_bb2_or_i17_i1866);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i1894_stall_local;
wire local_bb2_cmp77_i1894;

assign local_bb2_cmp77_i1894 = (local_bb2__33_i1879 > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u82_stall_local;
wire local_bb2_var__u82;

assign local_bb2_var__u82 = ($signed(local_bb2__33_i1879) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_cmp53_i1884_stall_local;
wire local_bb2_cmp53_i1884;

assign local_bb2_cmp53_i1884 = (local_bb2__37_i1883 > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp68_i1888_stall_local;
wire local_bb2_cmp68_i1888;

assign local_bb2_cmp68_i1888 = (local_bb2__37_i1883 < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i1890_stall_local;
wire [31:0] local_bb2_sub_i1890;

assign local_bb2_sub_i1890 = (local_bb2__37_i1883 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp71_not_i1905_stall_local;
wire local_bb2_cmp71_not_i1905;

assign local_bb2_cmp71_not_i1905 = (local_bb2__37_i1883 != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__35_i1332_stall_local;
wire [31:0] local_bb2__35_i1332;

assign local_bb2__35_i1332 = (local_bb2_tobool49_i1321 ? local_bb2__34_i1331 : local_bb2_or_i17_i1317);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i1345_stall_local;
wire local_bb2_cmp77_i1345;

assign local_bb2_cmp77_i1345 = (local_bb2__33_i1330 > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u83_stall_local;
wire local_bb2_var__u83;

assign local_bb2_var__u83 = ($signed(local_bb2__33_i1330) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2__35_i784_stall_local;
wire [31:0] local_bb2__35_i784;

assign local_bb2__35_i784 = (local_bb2_tobool49_i773 ? local_bb2__34_i783 : local_bb2_or_i17_i769);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i797_stall_local;
wire local_bb2_cmp77_i797;

assign local_bb2_cmp77_i797 = (local_bb2__33_i782 > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u84_stall_local;
wire local_bb2_var__u84;

assign local_bb2_var__u84 = ($signed(local_bb2__33_i782) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_cmp53_i787_stall_local;
wire local_bb2_cmp53_i787;

assign local_bb2_cmp53_i787 = (local_bb2__37_i786 > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp68_i791_stall_local;
wire local_bb2_cmp68_i791;

assign local_bb2_cmp68_i791 = (local_bb2__37_i786 < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i793_stall_local;
wire [31:0] local_bb2_sub_i793;

assign local_bb2_sub_i793 = (local_bb2__37_i786 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp71_not_i808_stall_local;
wire local_bb2_cmp71_not_i808;

assign local_bb2_cmp71_not_i808 = (local_bb2__37_i786 != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__35_i320_stall_local;
wire [31:0] local_bb2__35_i320;

assign local_bb2__35_i320 = (local_bb2_tobool49_i309 ? local_bb2__34_i319 : local_bb2_or_i17_i305);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i333_stall_local;
wire local_bb2_cmp77_i333;

assign local_bb2_cmp77_i333 = (local_bb2__33_i318 > 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u85_stall_local;
wire local_bb2_var__u85;

assign local_bb2_var__u85 = ($signed(local_bb2__33_i318) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i_stall_local;
wire [31:0] local_bb2_and75_i;

assign local_bb2_and75_i = (local_bb2__35_i & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and83_i_stall_local;
wire [31:0] local_bb2_and83_i;

assign local_bb2_and83_i = (local_bb2__35_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or581_i_stall_local;
wire local_bb2_or581_i;

assign local_bb2_or581_i = (rnode_168to169_bb2_var__u46_0_NO_SHIFT_REG | local_bb2_cmp53_i);

// This section implements an unregistered operation.
// 
wire local_bb2_and74_i_stall_local;
wire [31:0] local_bb2_and74_i;

assign local_bb2_and74_i = (local_bb2_sub_i + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i1432_stall_local;
wire [31:0] local_bb2_and75_i1432;

assign local_bb2_and75_i1432 = (local_bb2__35_i1424 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and83_i1438_stall_local;
wire [31:0] local_bb2_and83_i1438;

assign local_bb2_and83_i1438 = (local_bb2__35_i1424 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i884_stall_local;
wire [31:0] local_bb2_and75_i884;

assign local_bb2_and75_i884 = (local_bb2__35_i876 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and83_i890_stall_local;
wire [31:0] local_bb2_and83_i890;

assign local_bb2_and83_i890 = (local_bb2__35_i876 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i420_stall_local;
wire [31:0] local_bb2_and75_i420;

assign local_bb2_and75_i420 = (local_bb2__35_i412 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and83_i426_stall_local;
wire [31:0] local_bb2_and83_i426;

assign local_bb2_and83_i426 = (local_bb2__35_i412 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i1889_stall_local;
wire [31:0] local_bb2_and75_i1889;

assign local_bb2_and75_i1889 = (local_bb2__35_i1881 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and83_i1895_stall_local;
wire [31:0] local_bb2_and83_i1895;

assign local_bb2_and83_i1895 = (local_bb2__35_i1881 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or581_i1885_stall_local;
wire local_bb2_or581_i1885;

assign local_bb2_or581_i1885 = (rnode_168to169_bb2_var__u54_0_NO_SHIFT_REG | local_bb2_cmp53_i1884);

// This section implements an unregistered operation.
// 
wire local_bb2_and74_i1891_stall_local;
wire [31:0] local_bb2_and74_i1891;

assign local_bb2_and74_i1891 = (local_bb2_sub_i1890 + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i1340_stall_local;
wire [31:0] local_bb2_and75_i1340;

assign local_bb2_and75_i1340 = (local_bb2__35_i1332 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and83_i1346_stall_local;
wire [31:0] local_bb2_and83_i1346;

assign local_bb2_and83_i1346 = (local_bb2__35_i1332 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i792_stall_local;
wire [31:0] local_bb2_and75_i792;

assign local_bb2_and75_i792 = (local_bb2__35_i784 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and83_i798_stall_local;
wire [31:0] local_bb2_and83_i798;

assign local_bb2_and83_i798 = (local_bb2__35_i784 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or581_i788_stall_local;
wire local_bb2_or581_i788;

assign local_bb2_or581_i788 = (rnode_168to169_bb2_var__u58_0_NO_SHIFT_REG | local_bb2_cmp53_i787);

// This section implements an unregistered operation.
// 
wire local_bb2_and74_i794_stall_local;
wire [31:0] local_bb2_and74_i794;

assign local_bb2_and74_i794 = (local_bb2_sub_i793 + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i328_stall_local;
wire [31:0] local_bb2_and75_i328;

assign local_bb2_and75_i328 = (local_bb2__35_i320 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and83_i334_stall_local;
wire [31:0] local_bb2_and83_i334;

assign local_bb2_and83_i334 = (local_bb2__35_i320 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool84_i_stall_local;
wire local_bb2_tobool84_i;

assign local_bb2_tobool84_i = (local_bb2_and83_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool84_i1439_stall_local;
wire local_bb2_tobool84_i1439;

assign local_bb2_tobool84_i1439 = (local_bb2_and83_i1438 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool84_i891_stall_local;
wire local_bb2_tobool84_i891;

assign local_bb2_tobool84_i891 = (local_bb2_and83_i890 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool84_i427_stall_local;
wire local_bb2_tobool84_i427;

assign local_bb2_tobool84_i427 = (local_bb2_and83_i426 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool84_i1896_stall_local;
wire local_bb2_tobool84_i1896;

assign local_bb2_tobool84_i1896 = (local_bb2_and83_i1895 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool84_i1347_stall_local;
wire local_bb2_tobool84_i1347;

assign local_bb2_tobool84_i1347 = (local_bb2_and83_i1346 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool84_i799_stall_local;
wire local_bb2_tobool84_i799;

assign local_bb2_tobool84_i799 = (local_bb2_and83_i798 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool84_i335_stall_local;
wire local_bb2_tobool84_i335;

assign local_bb2_tobool84_i335 = (local_bb2_and83_i334 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i_valid_out;
wire local_bb2_cmp77_i_stall_in;
 reg local_bb2_cmp77_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp68_i_valid_out;
wire local_bb2_cmp68_i_stall_in;
 reg local_bb2_cmp68_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp71_not_i_valid_out;
wire local_bb2_cmp71_not_i_stall_in;
 reg local_bb2_cmp71_not_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_and75_i_valid_out;
wire local_bb2_and75_i_stall_in;
 reg local_bb2_and75_i_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i_valid_out;
wire local_bb2__39_i_stall_in;
 reg local_bb2__39_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_or581_i_valid_out;
wire local_bb2_or581_i_stall_in;
 reg local_bb2_or581_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_and74_i_valid_out;
wire local_bb2_and74_i_stall_in;
 reg local_bb2_and74_i_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i_inputs_ready;
wire local_bb2__39_i_stall_local;
wire local_bb2__39_i;

assign local_bb2__39_i_inputs_ready = (local_bb2_mul_i_i_valid_out_0_NO_SHIFT_REG & local_bb2_mul_i_i_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i_0_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i_0_valid_out_0_NO_SHIFT_REG & rnode_168to169_bb2_add_i_0_valid_out_2_NO_SHIFT_REG & rnode_168to169_bb2_var__u46_0_valid_out_NO_SHIFT_REG);
assign local_bb2__39_i = (local_bb2_tobool84_i & local_bb2_var__u78);
assign local_bb2_cmp77_i_valid_out = 1'b1;
assign local_bb2_cmp68_i_valid_out = 1'b1;
assign local_bb2_cmp71_not_i_valid_out = 1'b1;
assign local_bb2_and75_i_valid_out = 1'b1;
assign local_bb2__39_i_valid_out = 1'b1;
assign local_bb2_or581_i_valid_out = 1'b1;
assign local_bb2_and74_i_valid_out = 1'b1;
assign local_bb2_mul_i_i_stall_in_0 = 1'b0;
assign local_bb2_mul_i_i_stall_in_1 = 1'b0;
assign rnode_168to169_bb2_add_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u46_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp77_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp68_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp71_not_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and75_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__39_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_or581_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and74_i_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp77_i_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i_inputs_ready & (local_bb2_cmp77_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp77_i_stall_in)) & local_bb2__39_i_stall_local);
		local_bb2_cmp68_i_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i_inputs_ready & (local_bb2_cmp68_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp68_i_stall_in)) & local_bb2__39_i_stall_local);
		local_bb2_cmp71_not_i_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i_inputs_ready & (local_bb2_cmp71_not_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp71_not_i_stall_in)) & local_bb2__39_i_stall_local);
		local_bb2_and75_i_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i_inputs_ready & (local_bb2_and75_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_and75_i_stall_in)) & local_bb2__39_i_stall_local);
		local_bb2__39_i_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i_inputs_ready & (local_bb2__39_i_consumed_0_NO_SHIFT_REG | ~(local_bb2__39_i_stall_in)) & local_bb2__39_i_stall_local);
		local_bb2_or581_i_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i_inputs_ready & (local_bb2_or581_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_or581_i_stall_in)) & local_bb2__39_i_stall_local);
		local_bb2_and74_i_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i_inputs_ready & (local_bb2_and74_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_and74_i_stall_in)) & local_bb2__39_i_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i1437_valid_out;
wire local_bb2_cmp77_i1437_stall_in;
 reg local_bb2_cmp77_i1437_consumed_0_NO_SHIFT_REG;
wire local_bb2__37_i1426_valid_out;
wire local_bb2__37_i1426_stall_in;
 reg local_bb2__37_i1426_consumed_0_NO_SHIFT_REG;
wire local_bb2_and75_i1432_valid_out;
wire local_bb2_and75_i1432_stall_in;
 reg local_bb2_and75_i1432_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i1440_valid_out;
wire local_bb2__39_i1440_stall_in;
 reg local_bb2__39_i1440_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i1440_inputs_ready;
wire local_bb2__39_i1440_stall_local;
wire local_bb2__39_i1440;

assign local_bb2__39_i1440_inputs_ready = (local_bb2_mul_i_i1404_valid_out_0_NO_SHIFT_REG & local_bb2_mul_i_i1404_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i1411_0_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i1411_0_valid_out_0_NO_SHIFT_REG & rnode_168to169_bb2_add_i1411_0_valid_out_2_NO_SHIFT_REG);
assign local_bb2__39_i1440 = (local_bb2_tobool84_i1439 & local_bb2_var__u79);
assign local_bb2_cmp77_i1437_valid_out = 1'b1;
assign local_bb2__37_i1426_valid_out = 1'b1;
assign local_bb2_and75_i1432_valid_out = 1'b1;
assign local_bb2__39_i1440_valid_out = 1'b1;
assign local_bb2_mul_i_i1404_stall_in_0 = 1'b0;
assign local_bb2_mul_i_i1404_stall_in_1 = 1'b0;
assign rnode_168to169_bb2_add_i1411_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1411_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1411_0_stall_in_2_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp77_i1437_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__37_i1426_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and75_i1432_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__39_i1440_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp77_i1437_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1440_inputs_ready & (local_bb2_cmp77_i1437_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp77_i1437_stall_in)) & local_bb2__39_i1440_stall_local);
		local_bb2__37_i1426_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1440_inputs_ready & (local_bb2__37_i1426_consumed_0_NO_SHIFT_REG | ~(local_bb2__37_i1426_stall_in)) & local_bb2__39_i1440_stall_local);
		local_bb2_and75_i1432_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1440_inputs_ready & (local_bb2_and75_i1432_consumed_0_NO_SHIFT_REG | ~(local_bb2_and75_i1432_stall_in)) & local_bb2__39_i1440_stall_local);
		local_bb2__39_i1440_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1440_inputs_ready & (local_bb2__39_i1440_consumed_0_NO_SHIFT_REG | ~(local_bb2__39_i1440_stall_in)) & local_bb2__39_i1440_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i889_valid_out;
wire local_bb2_cmp77_i889_stall_in;
 reg local_bb2_cmp77_i889_consumed_0_NO_SHIFT_REG;
wire local_bb2__37_i878_valid_out;
wire local_bb2__37_i878_stall_in;
 reg local_bb2__37_i878_consumed_0_NO_SHIFT_REG;
wire local_bb2_and75_i884_valid_out;
wire local_bb2_and75_i884_stall_in;
 reg local_bb2_and75_i884_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i892_valid_out;
wire local_bb2__39_i892_stall_in;
 reg local_bb2__39_i892_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i892_inputs_ready;
wire local_bb2__39_i892_stall_local;
wire local_bb2__39_i892;

assign local_bb2__39_i892_inputs_ready = (local_bb2_mul_i_i856_valid_out_0_NO_SHIFT_REG & local_bb2_mul_i_i856_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i863_0_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i863_0_valid_out_0_NO_SHIFT_REG & rnode_168to169_bb2_add_i863_0_valid_out_2_NO_SHIFT_REG);
assign local_bb2__39_i892 = (local_bb2_tobool84_i891 & local_bb2_var__u80);
assign local_bb2_cmp77_i889_valid_out = 1'b1;
assign local_bb2__37_i878_valid_out = 1'b1;
assign local_bb2_and75_i884_valid_out = 1'b1;
assign local_bb2__39_i892_valid_out = 1'b1;
assign local_bb2_mul_i_i856_stall_in_0 = 1'b0;
assign local_bb2_mul_i_i856_stall_in_1 = 1'b0;
assign rnode_168to169_bb2_add_i863_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i863_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i863_0_stall_in_2_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp77_i889_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__37_i878_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and75_i884_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__39_i892_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp77_i889_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i892_inputs_ready & (local_bb2_cmp77_i889_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp77_i889_stall_in)) & local_bb2__39_i892_stall_local);
		local_bb2__37_i878_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i892_inputs_ready & (local_bb2__37_i878_consumed_0_NO_SHIFT_REG | ~(local_bb2__37_i878_stall_in)) & local_bb2__39_i892_stall_local);
		local_bb2_and75_i884_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i892_inputs_ready & (local_bb2_and75_i884_consumed_0_NO_SHIFT_REG | ~(local_bb2_and75_i884_stall_in)) & local_bb2__39_i892_stall_local);
		local_bb2__39_i892_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i892_inputs_ready & (local_bb2__39_i892_consumed_0_NO_SHIFT_REG | ~(local_bb2__39_i892_stall_in)) & local_bb2__39_i892_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i425_valid_out;
wire local_bb2_cmp77_i425_stall_in;
 reg local_bb2_cmp77_i425_consumed_0_NO_SHIFT_REG;
wire local_bb2__37_i414_valid_out;
wire local_bb2__37_i414_stall_in;
 reg local_bb2__37_i414_consumed_0_NO_SHIFT_REG;
wire local_bb2_and75_i420_valid_out;
wire local_bb2_and75_i420_stall_in;
 reg local_bb2_and75_i420_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i428_valid_out;
wire local_bb2__39_i428_stall_in;
 reg local_bb2__39_i428_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i428_inputs_ready;
wire local_bb2__39_i428_stall_local;
wire local_bb2__39_i428;

assign local_bb2__39_i428_inputs_ready = (local_bb2_mul_i_i392_valid_out_0_NO_SHIFT_REG & local_bb2_mul_i_i392_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i399_0_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i399_0_valid_out_0_NO_SHIFT_REG & rnode_168to169_bb2_add_i399_0_valid_out_2_NO_SHIFT_REG);
assign local_bb2__39_i428 = (local_bb2_tobool84_i427 & local_bb2_var__u81);
assign local_bb2_cmp77_i425_valid_out = 1'b1;
assign local_bb2__37_i414_valid_out = 1'b1;
assign local_bb2_and75_i420_valid_out = 1'b1;
assign local_bb2__39_i428_valid_out = 1'b1;
assign local_bb2_mul_i_i392_stall_in_0 = 1'b0;
assign local_bb2_mul_i_i392_stall_in_1 = 1'b0;
assign rnode_168to169_bb2_add_i399_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i399_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i399_0_stall_in_2_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp77_i425_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__37_i414_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and75_i420_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__39_i428_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp77_i425_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i428_inputs_ready & (local_bb2_cmp77_i425_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp77_i425_stall_in)) & local_bb2__39_i428_stall_local);
		local_bb2__37_i414_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i428_inputs_ready & (local_bb2__37_i414_consumed_0_NO_SHIFT_REG | ~(local_bb2__37_i414_stall_in)) & local_bb2__39_i428_stall_local);
		local_bb2_and75_i420_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i428_inputs_ready & (local_bb2_and75_i420_consumed_0_NO_SHIFT_REG | ~(local_bb2_and75_i420_stall_in)) & local_bb2__39_i428_stall_local);
		local_bb2__39_i428_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i428_inputs_ready & (local_bb2__39_i428_consumed_0_NO_SHIFT_REG | ~(local_bb2__39_i428_stall_in)) & local_bb2__39_i428_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i1894_valid_out;
wire local_bb2_cmp77_i1894_stall_in;
 reg local_bb2_cmp77_i1894_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp68_i1888_valid_out;
wire local_bb2_cmp68_i1888_stall_in;
 reg local_bb2_cmp68_i1888_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp71_not_i1905_valid_out;
wire local_bb2_cmp71_not_i1905_stall_in;
 reg local_bb2_cmp71_not_i1905_consumed_0_NO_SHIFT_REG;
wire local_bb2_and75_i1889_valid_out;
wire local_bb2_and75_i1889_stall_in;
 reg local_bb2_and75_i1889_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i1897_valid_out;
wire local_bb2__39_i1897_stall_in;
 reg local_bb2__39_i1897_consumed_0_NO_SHIFT_REG;
wire local_bb2_or581_i1885_valid_out;
wire local_bb2_or581_i1885_stall_in;
 reg local_bb2_or581_i1885_consumed_0_NO_SHIFT_REG;
wire local_bb2_and74_i1891_valid_out;
wire local_bb2_and74_i1891_stall_in;
 reg local_bb2_and74_i1891_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i1897_inputs_ready;
wire local_bb2__39_i1897_stall_local;
wire local_bb2__39_i1897;

assign local_bb2__39_i1897_inputs_ready = (local_bb2_mul_i_i1861_valid_out_0_NO_SHIFT_REG & local_bb2_mul_i_i1861_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i1868_0_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i1868_0_valid_out_0_NO_SHIFT_REG & rnode_168to169_bb2_add_i1868_0_valid_out_2_NO_SHIFT_REG & rnode_168to169_bb2_var__u54_0_valid_out_NO_SHIFT_REG);
assign local_bb2__39_i1897 = (local_bb2_tobool84_i1896 & local_bb2_var__u82);
assign local_bb2_cmp77_i1894_valid_out = 1'b1;
assign local_bb2_cmp68_i1888_valid_out = 1'b1;
assign local_bb2_cmp71_not_i1905_valid_out = 1'b1;
assign local_bb2_and75_i1889_valid_out = 1'b1;
assign local_bb2__39_i1897_valid_out = 1'b1;
assign local_bb2_or581_i1885_valid_out = 1'b1;
assign local_bb2_and74_i1891_valid_out = 1'b1;
assign local_bb2_mul_i_i1861_stall_in_0 = 1'b0;
assign local_bb2_mul_i_i1861_stall_in_1 = 1'b0;
assign rnode_168to169_bb2_add_i1868_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1868_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1868_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u54_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp77_i1894_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp68_i1888_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp71_not_i1905_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and75_i1889_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__39_i1897_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_or581_i1885_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and74_i1891_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp77_i1894_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1897_inputs_ready & (local_bb2_cmp77_i1894_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp77_i1894_stall_in)) & local_bb2__39_i1897_stall_local);
		local_bb2_cmp68_i1888_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1897_inputs_ready & (local_bb2_cmp68_i1888_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp68_i1888_stall_in)) & local_bb2__39_i1897_stall_local);
		local_bb2_cmp71_not_i1905_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1897_inputs_ready & (local_bb2_cmp71_not_i1905_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp71_not_i1905_stall_in)) & local_bb2__39_i1897_stall_local);
		local_bb2_and75_i1889_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1897_inputs_ready & (local_bb2_and75_i1889_consumed_0_NO_SHIFT_REG | ~(local_bb2_and75_i1889_stall_in)) & local_bb2__39_i1897_stall_local);
		local_bb2__39_i1897_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1897_inputs_ready & (local_bb2__39_i1897_consumed_0_NO_SHIFT_REG | ~(local_bb2__39_i1897_stall_in)) & local_bb2__39_i1897_stall_local);
		local_bb2_or581_i1885_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1897_inputs_ready & (local_bb2_or581_i1885_consumed_0_NO_SHIFT_REG | ~(local_bb2_or581_i1885_stall_in)) & local_bb2__39_i1897_stall_local);
		local_bb2_and74_i1891_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1897_inputs_ready & (local_bb2_and74_i1891_consumed_0_NO_SHIFT_REG | ~(local_bb2_and74_i1891_stall_in)) & local_bb2__39_i1897_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i1345_valid_out;
wire local_bb2_cmp77_i1345_stall_in;
 reg local_bb2_cmp77_i1345_consumed_0_NO_SHIFT_REG;
wire local_bb2__37_i1334_valid_out;
wire local_bb2__37_i1334_stall_in;
 reg local_bb2__37_i1334_consumed_0_NO_SHIFT_REG;
wire local_bb2_and75_i1340_valid_out;
wire local_bb2_and75_i1340_stall_in;
 reg local_bb2_and75_i1340_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i1348_valid_out;
wire local_bb2__39_i1348_stall_in;
 reg local_bb2__39_i1348_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i1348_inputs_ready;
wire local_bb2__39_i1348_stall_local;
wire local_bb2__39_i1348;

assign local_bb2__39_i1348_inputs_ready = (local_bb2_mul_i_i1312_valid_out_0_NO_SHIFT_REG & local_bb2_mul_i_i1312_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i1319_0_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i1319_0_valid_out_0_NO_SHIFT_REG & rnode_168to169_bb2_add_i1319_0_valid_out_2_NO_SHIFT_REG);
assign local_bb2__39_i1348 = (local_bb2_tobool84_i1347 & local_bb2_var__u83);
assign local_bb2_cmp77_i1345_valid_out = 1'b1;
assign local_bb2__37_i1334_valid_out = 1'b1;
assign local_bb2_and75_i1340_valid_out = 1'b1;
assign local_bb2__39_i1348_valid_out = 1'b1;
assign local_bb2_mul_i_i1312_stall_in_0 = 1'b0;
assign local_bb2_mul_i_i1312_stall_in_1 = 1'b0;
assign rnode_168to169_bb2_add_i1319_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1319_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i1319_0_stall_in_2_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp77_i1345_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__37_i1334_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and75_i1340_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__39_i1348_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp77_i1345_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1348_inputs_ready & (local_bb2_cmp77_i1345_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp77_i1345_stall_in)) & local_bb2__39_i1348_stall_local);
		local_bb2__37_i1334_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1348_inputs_ready & (local_bb2__37_i1334_consumed_0_NO_SHIFT_REG | ~(local_bb2__37_i1334_stall_in)) & local_bb2__39_i1348_stall_local);
		local_bb2_and75_i1340_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1348_inputs_ready & (local_bb2_and75_i1340_consumed_0_NO_SHIFT_REG | ~(local_bb2_and75_i1340_stall_in)) & local_bb2__39_i1348_stall_local);
		local_bb2__39_i1348_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i1348_inputs_ready & (local_bb2__39_i1348_consumed_0_NO_SHIFT_REG | ~(local_bb2__39_i1348_stall_in)) & local_bb2__39_i1348_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i797_valid_out;
wire local_bb2_cmp77_i797_stall_in;
 reg local_bb2_cmp77_i797_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp68_i791_valid_out;
wire local_bb2_cmp68_i791_stall_in;
 reg local_bb2_cmp68_i791_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp71_not_i808_valid_out;
wire local_bb2_cmp71_not_i808_stall_in;
 reg local_bb2_cmp71_not_i808_consumed_0_NO_SHIFT_REG;
wire local_bb2_and75_i792_valid_out;
wire local_bb2_and75_i792_stall_in;
 reg local_bb2_and75_i792_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i800_valid_out;
wire local_bb2__39_i800_stall_in;
 reg local_bb2__39_i800_consumed_0_NO_SHIFT_REG;
wire local_bb2_or581_i788_valid_out;
wire local_bb2_or581_i788_stall_in;
 reg local_bb2_or581_i788_consumed_0_NO_SHIFT_REG;
wire local_bb2_and74_i794_valid_out;
wire local_bb2_and74_i794_stall_in;
 reg local_bb2_and74_i794_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i800_inputs_ready;
wire local_bb2__39_i800_stall_local;
wire local_bb2__39_i800;

assign local_bb2__39_i800_inputs_ready = (local_bb2_mul_i_i764_valid_out_0_NO_SHIFT_REG & local_bb2_mul_i_i764_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i771_0_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i771_0_valid_out_0_NO_SHIFT_REG & rnode_168to169_bb2_add_i771_0_valid_out_2_NO_SHIFT_REG & rnode_168to169_bb2_var__u58_0_valid_out_NO_SHIFT_REG);
assign local_bb2__39_i800 = (local_bb2_tobool84_i799 & local_bb2_var__u84);
assign local_bb2_cmp77_i797_valid_out = 1'b1;
assign local_bb2_cmp68_i791_valid_out = 1'b1;
assign local_bb2_cmp71_not_i808_valid_out = 1'b1;
assign local_bb2_and75_i792_valid_out = 1'b1;
assign local_bb2__39_i800_valid_out = 1'b1;
assign local_bb2_or581_i788_valid_out = 1'b1;
assign local_bb2_and74_i794_valid_out = 1'b1;
assign local_bb2_mul_i_i764_stall_in_0 = 1'b0;
assign local_bb2_mul_i_i764_stall_in_1 = 1'b0;
assign rnode_168to169_bb2_add_i771_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i771_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i771_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_var__u58_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp77_i797_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp68_i791_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp71_not_i808_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and75_i792_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__39_i800_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_or581_i788_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and74_i794_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp77_i797_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i800_inputs_ready & (local_bb2_cmp77_i797_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp77_i797_stall_in)) & local_bb2__39_i800_stall_local);
		local_bb2_cmp68_i791_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i800_inputs_ready & (local_bb2_cmp68_i791_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp68_i791_stall_in)) & local_bb2__39_i800_stall_local);
		local_bb2_cmp71_not_i808_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i800_inputs_ready & (local_bb2_cmp71_not_i808_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp71_not_i808_stall_in)) & local_bb2__39_i800_stall_local);
		local_bb2_and75_i792_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i800_inputs_ready & (local_bb2_and75_i792_consumed_0_NO_SHIFT_REG | ~(local_bb2_and75_i792_stall_in)) & local_bb2__39_i800_stall_local);
		local_bb2__39_i800_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i800_inputs_ready & (local_bb2__39_i800_consumed_0_NO_SHIFT_REG | ~(local_bb2__39_i800_stall_in)) & local_bb2__39_i800_stall_local);
		local_bb2_or581_i788_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i800_inputs_ready & (local_bb2_or581_i788_consumed_0_NO_SHIFT_REG | ~(local_bb2_or581_i788_stall_in)) & local_bb2__39_i800_stall_local);
		local_bb2_and74_i794_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i800_inputs_ready & (local_bb2_and74_i794_consumed_0_NO_SHIFT_REG | ~(local_bb2_and74_i794_stall_in)) & local_bb2__39_i800_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i333_valid_out;
wire local_bb2_cmp77_i333_stall_in;
 reg local_bb2_cmp77_i333_consumed_0_NO_SHIFT_REG;
wire local_bb2__37_i322_valid_out;
wire local_bb2__37_i322_stall_in;
 reg local_bb2__37_i322_consumed_0_NO_SHIFT_REG;
wire local_bb2_and75_i328_valid_out;
wire local_bb2_and75_i328_stall_in;
 reg local_bb2_and75_i328_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i336_valid_out;
wire local_bb2__39_i336_stall_in;
 reg local_bb2__39_i336_consumed_0_NO_SHIFT_REG;
wire local_bb2__39_i336_inputs_ready;
wire local_bb2__39_i336_stall_local;
wire local_bb2__39_i336;

assign local_bb2__39_i336_inputs_ready = (local_bb2_mul_i_i300_valid_out_0_NO_SHIFT_REG & local_bb2_mul_i_i300_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i307_0_valid_out_1_NO_SHIFT_REG & rnode_168to169_bb2_add_i307_0_valid_out_0_NO_SHIFT_REG & rnode_168to169_bb2_add_i307_0_valid_out_2_NO_SHIFT_REG);
assign local_bb2__39_i336 = (local_bb2_tobool84_i335 & local_bb2_var__u85);
assign local_bb2_cmp77_i333_valid_out = 1'b1;
assign local_bb2__37_i322_valid_out = 1'b1;
assign local_bb2_and75_i328_valid_out = 1'b1;
assign local_bb2__39_i336_valid_out = 1'b1;
assign local_bb2_mul_i_i300_stall_in_0 = 1'b0;
assign local_bb2_mul_i_i300_stall_in_1 = 1'b0;
assign rnode_168to169_bb2_add_i307_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i307_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_168to169_bb2_add_i307_0_stall_in_2_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp77_i333_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__37_i322_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and75_i328_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__39_i336_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp77_i333_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i336_inputs_ready & (local_bb2_cmp77_i333_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp77_i333_stall_in)) & local_bb2__39_i336_stall_local);
		local_bb2__37_i322_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i336_inputs_ready & (local_bb2__37_i322_consumed_0_NO_SHIFT_REG | ~(local_bb2__37_i322_stall_in)) & local_bb2__39_i336_stall_local);
		local_bb2_and75_i328_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i336_inputs_ready & (local_bb2_and75_i328_consumed_0_NO_SHIFT_REG | ~(local_bb2_and75_i328_stall_in)) & local_bb2__39_i336_stall_local);
		local_bb2__39_i336_consumed_0_NO_SHIFT_REG <= (local_bb2__39_i336_inputs_ready & (local_bb2__39_i336_consumed_0_NO_SHIFT_REG | ~(local_bb2__39_i336_stall_in)) & local_bb2__39_i336_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp77_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp77_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp77_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp77_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp77_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp77_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp77_i),
	.data_out(rnode_169to170_bb2_cmp77_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp77_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp77_i_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp77_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp77_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp77_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp77_i_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp77_i_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp77_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp77_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp68_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp68_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp68_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp68_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp68_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp68_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp68_i),
	.data_out(rnode_169to170_bb2_cmp68_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp68_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp68_i_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp68_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp68_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp68_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp68_i_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp68_i_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp68_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp68_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp68_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp71_not_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp71_not_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp71_not_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp71_not_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp71_not_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp71_not_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp71_not_i),
	.data_out(rnode_169to170_bb2_cmp71_not_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp71_not_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp71_not_i_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp71_not_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp71_not_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp71_not_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp71_not_i_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp71_not_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp71_not_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and75_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and75_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and75_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and75_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and75_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and75_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and75_i),
	.data_out(rnode_169to170_bb2_and75_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and75_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and75_i_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and75_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and75_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and75_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and75_i_stall_in = 1'b0;
assign rnode_169to170_bb2_and75_i_0_NO_SHIFT_REG = rnode_169to170_bb2_and75_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and75_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__39_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__39_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__39_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__39_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__39_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__39_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__39_i),
	.data_out(rnode_169to170_bb2__39_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__39_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__39_i_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__39_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__39_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__39_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__39_i_stall_in = 1'b0;
assign rnode_169to170_bb2__39_i_0_NO_SHIFT_REG = rnode_169to170_bb2__39_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__39_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_or581_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_valid_out_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_stall_in_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_or581_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_or581_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_or581_i_0_stall_in_0_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_or581_i_0_valid_out_0_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_or581_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_or581_i),
	.data_out(rnode_169to170_bb2_or581_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_or581_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_or581_i_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_or581_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_or581_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_or581_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or581_i_stall_in = 1'b0;
assign rnode_169to170_bb2_or581_i_0_stall_in_0_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2_or581_i_0_NO_SHIFT_REG = rnode_169to170_bb2_or581_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_or581_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2_or581_i_1_NO_SHIFT_REG = rnode_169to170_bb2_or581_i_0_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and74_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and74_i_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and74_i_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and74_i_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and74_i_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and74_i_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and74_i_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and74_i_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and74_i),
	.data_out(rnode_169to170_bb2_and74_i_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and74_i_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and74_i_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and74_i_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and74_i_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and74_i_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and74_i_stall_in = 1'b0;
assign rnode_169to170_bb2_and74_i_0_NO_SHIFT_REG = rnode_169to170_bb2_and74_i_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and74_i_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and74_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp77_i1437_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1437_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1437_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1437_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1437_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1437_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1437_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1437_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp77_i1437_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp77_i1437_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp77_i1437_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp77_i1437_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp77_i1437_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp77_i1437),
	.data_out(rnode_169to170_bb2_cmp77_i1437_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp77_i1437_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp77_i1437_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp77_i1437_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp77_i1437_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp77_i1437_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp77_i1437_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp77_i1437_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp77_i1437_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp77_i1437_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i1437_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__37_i1426_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1426_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1426_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1426_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1426_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1426_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_valid_out_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_stall_in_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1426_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__37_i1426_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__37_i1426_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__37_i1426_0_stall_in_0_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__37_i1426_0_valid_out_0_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__37_i1426_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__37_i1426),
	.data_out(rnode_169to170_bb2__37_i1426_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__37_i1426_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__37_i1426_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2__37_i1426_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__37_i1426_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__37_i1426_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__37_i1426_stall_in = 1'b0;
assign rnode_169to170_bb2__37_i1426_0_stall_in_0_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1426_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i1426_0_NO_SHIFT_REG = rnode_169to170_bb2__37_i1426_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i1426_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i1426_1_NO_SHIFT_REG = rnode_169to170_bb2__37_i1426_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i1426_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i1426_2_NO_SHIFT_REG = rnode_169to170_bb2__37_i1426_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i1426_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i1426_3_NO_SHIFT_REG = rnode_169to170_bb2__37_i1426_0_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and75_i1432_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1432_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i1432_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1432_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i1432_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1432_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1432_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1432_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and75_i1432_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and75_i1432_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and75_i1432_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and75_i1432_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and75_i1432_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and75_i1432),
	.data_out(rnode_169to170_bb2_and75_i1432_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and75_i1432_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and75_i1432_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and75_i1432_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and75_i1432_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and75_i1432_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and75_i1432_stall_in = 1'b0;
assign rnode_169to170_bb2_and75_i1432_0_NO_SHIFT_REG = rnode_169to170_bb2_and75_i1432_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and75_i1432_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i1432_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__39_i1440_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1440_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1440_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1440_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1440_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1440_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1440_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1440_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__39_i1440_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__39_i1440_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__39_i1440_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__39_i1440_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__39_i1440_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__39_i1440),
	.data_out(rnode_169to170_bb2__39_i1440_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__39_i1440_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__39_i1440_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__39_i1440_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__39_i1440_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__39_i1440_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__39_i1440_stall_in = 1'b0;
assign rnode_169to170_bb2__39_i1440_0_NO_SHIFT_REG = rnode_169to170_bb2__39_i1440_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__39_i1440_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i1440_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp77_i889_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i889_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i889_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i889_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i889_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i889_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i889_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i889_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp77_i889_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp77_i889_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp77_i889_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp77_i889_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp77_i889_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp77_i889),
	.data_out(rnode_169to170_bb2_cmp77_i889_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp77_i889_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp77_i889_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp77_i889_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp77_i889_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp77_i889_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp77_i889_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp77_i889_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp77_i889_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp77_i889_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i889_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__37_i878_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i878_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i878_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i878_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i878_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i878_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_valid_out_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_stall_in_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i878_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__37_i878_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__37_i878_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__37_i878_0_stall_in_0_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__37_i878_0_valid_out_0_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__37_i878_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__37_i878),
	.data_out(rnode_169to170_bb2__37_i878_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__37_i878_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__37_i878_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2__37_i878_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__37_i878_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__37_i878_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__37_i878_stall_in = 1'b0;
assign rnode_169to170_bb2__37_i878_0_stall_in_0_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i878_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i878_0_NO_SHIFT_REG = rnode_169to170_bb2__37_i878_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i878_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i878_1_NO_SHIFT_REG = rnode_169to170_bb2__37_i878_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i878_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i878_2_NO_SHIFT_REG = rnode_169to170_bb2__37_i878_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i878_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i878_3_NO_SHIFT_REG = rnode_169to170_bb2__37_i878_0_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and75_i884_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i884_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i884_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i884_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i884_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i884_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i884_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i884_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and75_i884_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and75_i884_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and75_i884_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and75_i884_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and75_i884_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and75_i884),
	.data_out(rnode_169to170_bb2_and75_i884_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and75_i884_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and75_i884_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and75_i884_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and75_i884_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and75_i884_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and75_i884_stall_in = 1'b0;
assign rnode_169to170_bb2_and75_i884_0_NO_SHIFT_REG = rnode_169to170_bb2_and75_i884_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and75_i884_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i884_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__39_i892_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i892_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i892_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i892_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i892_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i892_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i892_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i892_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__39_i892_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__39_i892_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__39_i892_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__39_i892_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__39_i892_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__39_i892),
	.data_out(rnode_169to170_bb2__39_i892_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__39_i892_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__39_i892_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__39_i892_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__39_i892_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__39_i892_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__39_i892_stall_in = 1'b0;
assign rnode_169to170_bb2__39_i892_0_NO_SHIFT_REG = rnode_169to170_bb2__39_i892_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__39_i892_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i892_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp77_i425_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i425_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i425_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i425_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i425_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i425_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i425_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i425_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp77_i425_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp77_i425_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp77_i425_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp77_i425_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp77_i425_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp77_i425),
	.data_out(rnode_169to170_bb2_cmp77_i425_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp77_i425_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp77_i425_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp77_i425_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp77_i425_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp77_i425_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp77_i425_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp77_i425_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp77_i425_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp77_i425_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i425_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__37_i414_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i414_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i414_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i414_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i414_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i414_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_valid_out_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_stall_in_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i414_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__37_i414_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__37_i414_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__37_i414_0_stall_in_0_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__37_i414_0_valid_out_0_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__37_i414_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__37_i414),
	.data_out(rnode_169to170_bb2__37_i414_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__37_i414_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__37_i414_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2__37_i414_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__37_i414_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__37_i414_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__37_i414_stall_in = 1'b0;
assign rnode_169to170_bb2__37_i414_0_stall_in_0_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i414_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i414_0_NO_SHIFT_REG = rnode_169to170_bb2__37_i414_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i414_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i414_1_NO_SHIFT_REG = rnode_169to170_bb2__37_i414_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i414_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i414_2_NO_SHIFT_REG = rnode_169to170_bb2__37_i414_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i414_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i414_3_NO_SHIFT_REG = rnode_169to170_bb2__37_i414_0_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and75_i420_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i420_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i420_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i420_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i420_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i420_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i420_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i420_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and75_i420_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and75_i420_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and75_i420_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and75_i420_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and75_i420_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and75_i420),
	.data_out(rnode_169to170_bb2_and75_i420_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and75_i420_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and75_i420_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and75_i420_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and75_i420_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and75_i420_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and75_i420_stall_in = 1'b0;
assign rnode_169to170_bb2_and75_i420_0_NO_SHIFT_REG = rnode_169to170_bb2_and75_i420_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and75_i420_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i420_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__39_i428_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i428_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i428_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i428_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i428_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i428_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i428_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i428_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__39_i428_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__39_i428_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__39_i428_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__39_i428_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__39_i428_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__39_i428),
	.data_out(rnode_169to170_bb2__39_i428_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__39_i428_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__39_i428_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__39_i428_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__39_i428_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__39_i428_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__39_i428_stall_in = 1'b0;
assign rnode_169to170_bb2__39_i428_0_NO_SHIFT_REG = rnode_169to170_bb2__39_i428_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__39_i428_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i428_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp77_i1894_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1894_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1894_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1894_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1894_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1894_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1894_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1894_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp77_i1894_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp77_i1894_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp77_i1894_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp77_i1894_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp77_i1894_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp77_i1894),
	.data_out(rnode_169to170_bb2_cmp77_i1894_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp77_i1894_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp77_i1894_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp77_i1894_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp77_i1894_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp77_i1894_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp77_i1894_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp77_i1894_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp77_i1894_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp77_i1894_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i1894_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp68_i1888_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i1888_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i1888_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i1888_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i1888_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i1888_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i1888_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i1888_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp68_i1888_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp68_i1888_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp68_i1888_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp68_i1888_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp68_i1888_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp68_i1888),
	.data_out(rnode_169to170_bb2_cmp68_i1888_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp68_i1888_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp68_i1888_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp68_i1888_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp68_i1888_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp68_i1888_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp68_i1888_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp68_i1888_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp68_i1888_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp68_i1888_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp68_i1888_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp71_not_i1905_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i1905_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i1905_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i1905_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i1905_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i1905_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp71_not_i1905_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp71_not_i1905_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp71_not_i1905_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp71_not_i1905),
	.data_out(rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp71_not_i1905_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i1905_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp71_not_i1905_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp71_not_i1905_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i1905_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and75_i1889_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1889_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i1889_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1889_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i1889_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1889_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1889_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1889_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and75_i1889_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and75_i1889_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and75_i1889_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and75_i1889_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and75_i1889_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and75_i1889),
	.data_out(rnode_169to170_bb2_and75_i1889_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and75_i1889_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and75_i1889_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and75_i1889_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and75_i1889_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and75_i1889_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and75_i1889_stall_in = 1'b0;
assign rnode_169to170_bb2_and75_i1889_0_NO_SHIFT_REG = rnode_169to170_bb2_and75_i1889_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and75_i1889_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i1889_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__39_i1897_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1897_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1897_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1897_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1897_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1897_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1897_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1897_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__39_i1897_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__39_i1897_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__39_i1897_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__39_i1897_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__39_i1897_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__39_i1897),
	.data_out(rnode_169to170_bb2__39_i1897_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__39_i1897_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__39_i1897_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__39_i1897_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__39_i1897_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__39_i1897_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__39_i1897_stall_in = 1'b0;
assign rnode_169to170_bb2__39_i1897_0_NO_SHIFT_REG = rnode_169to170_bb2__39_i1897_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__39_i1897_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i1897_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_or581_i1885_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_valid_out_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_stall_in_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i1885_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_or581_i1885_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_or581_i1885_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_or581_i1885_0_stall_in_0_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_or581_i1885_0_valid_out_0_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_or581_i1885_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_or581_i1885),
	.data_out(rnode_169to170_bb2_or581_i1885_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_or581_i1885_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_or581_i1885_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_or581_i1885_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_or581_i1885_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_or581_i1885_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or581_i1885_stall_in = 1'b0;
assign rnode_169to170_bb2_or581_i1885_0_stall_in_0_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i1885_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2_or581_i1885_0_NO_SHIFT_REG = rnode_169to170_bb2_or581_i1885_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_or581_i1885_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2_or581_i1885_1_NO_SHIFT_REG = rnode_169to170_bb2_or581_i1885_0_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and74_i1891_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i1891_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and74_i1891_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i1891_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and74_i1891_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i1891_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i1891_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i1891_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and74_i1891_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and74_i1891_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and74_i1891_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and74_i1891_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and74_i1891_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and74_i1891),
	.data_out(rnode_169to170_bb2_and74_i1891_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and74_i1891_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and74_i1891_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and74_i1891_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and74_i1891_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and74_i1891_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and74_i1891_stall_in = 1'b0;
assign rnode_169to170_bb2_and74_i1891_0_NO_SHIFT_REG = rnode_169to170_bb2_and74_i1891_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and74_i1891_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and74_i1891_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp77_i1345_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1345_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1345_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1345_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1345_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1345_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1345_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i1345_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp77_i1345_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp77_i1345_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp77_i1345_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp77_i1345_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp77_i1345_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp77_i1345),
	.data_out(rnode_169to170_bb2_cmp77_i1345_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp77_i1345_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp77_i1345_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp77_i1345_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp77_i1345_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp77_i1345_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp77_i1345_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp77_i1345_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp77_i1345_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp77_i1345_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i1345_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__37_i1334_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1334_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1334_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1334_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1334_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i1334_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_valid_out_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_stall_in_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i1334_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__37_i1334_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__37_i1334_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__37_i1334_0_stall_in_0_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__37_i1334_0_valid_out_0_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__37_i1334_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__37_i1334),
	.data_out(rnode_169to170_bb2__37_i1334_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__37_i1334_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__37_i1334_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2__37_i1334_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__37_i1334_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__37_i1334_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__37_i1334_stall_in = 1'b0;
assign rnode_169to170_bb2__37_i1334_0_stall_in_0_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1334_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i1334_0_NO_SHIFT_REG = rnode_169to170_bb2__37_i1334_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i1334_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i1334_1_NO_SHIFT_REG = rnode_169to170_bb2__37_i1334_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i1334_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i1334_2_NO_SHIFT_REG = rnode_169to170_bb2__37_i1334_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i1334_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i1334_3_NO_SHIFT_REG = rnode_169to170_bb2__37_i1334_0_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and75_i1340_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1340_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i1340_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1340_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i1340_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1340_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1340_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i1340_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and75_i1340_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and75_i1340_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and75_i1340_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and75_i1340_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and75_i1340_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and75_i1340),
	.data_out(rnode_169to170_bb2_and75_i1340_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and75_i1340_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and75_i1340_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and75_i1340_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and75_i1340_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and75_i1340_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and75_i1340_stall_in = 1'b0;
assign rnode_169to170_bb2_and75_i1340_0_NO_SHIFT_REG = rnode_169to170_bb2_and75_i1340_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and75_i1340_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i1340_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__39_i1348_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1348_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1348_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1348_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1348_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1348_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1348_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i1348_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__39_i1348_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__39_i1348_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__39_i1348_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__39_i1348_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__39_i1348_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__39_i1348),
	.data_out(rnode_169to170_bb2__39_i1348_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__39_i1348_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__39_i1348_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__39_i1348_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__39_i1348_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__39_i1348_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__39_i1348_stall_in = 1'b0;
assign rnode_169to170_bb2__39_i1348_0_NO_SHIFT_REG = rnode_169to170_bb2__39_i1348_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__39_i1348_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i1348_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp77_i797_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i797_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i797_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i797_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i797_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i797_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i797_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i797_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp77_i797_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp77_i797_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp77_i797_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp77_i797_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp77_i797_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp77_i797),
	.data_out(rnode_169to170_bb2_cmp77_i797_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp77_i797_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp77_i797_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp77_i797_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp77_i797_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp77_i797_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp77_i797_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp77_i797_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp77_i797_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp77_i797_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i797_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp68_i791_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i791_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i791_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i791_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i791_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i791_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i791_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp68_i791_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp68_i791_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp68_i791_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp68_i791_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp68_i791_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp68_i791_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp68_i791),
	.data_out(rnode_169to170_bb2_cmp68_i791_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp68_i791_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp68_i791_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp68_i791_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp68_i791_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp68_i791_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp68_i791_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp68_i791_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp68_i791_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp68_i791_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp68_i791_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp71_not_i808_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i808_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i808_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i808_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i808_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i808_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i808_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp71_not_i808_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp71_not_i808_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp71_not_i808_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp71_not_i808_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp71_not_i808_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp71_not_i808_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp71_not_i808),
	.data_out(rnode_169to170_bb2_cmp71_not_i808_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp71_not_i808_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp71_not_i808_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp71_not_i808_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp71_not_i808_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp71_not_i808_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp71_not_i808_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i808_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp71_not_i808_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp71_not_i808_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i808_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and75_i792_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i792_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i792_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i792_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i792_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i792_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i792_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i792_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and75_i792_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and75_i792_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and75_i792_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and75_i792_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and75_i792_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and75_i792),
	.data_out(rnode_169to170_bb2_and75_i792_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and75_i792_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and75_i792_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and75_i792_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and75_i792_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and75_i792_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and75_i792_stall_in = 1'b0;
assign rnode_169to170_bb2_and75_i792_0_NO_SHIFT_REG = rnode_169to170_bb2_and75_i792_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and75_i792_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i792_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__39_i800_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i800_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i800_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i800_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i800_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i800_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i800_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i800_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__39_i800_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__39_i800_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__39_i800_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__39_i800_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__39_i800_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__39_i800),
	.data_out(rnode_169to170_bb2__39_i800_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__39_i800_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__39_i800_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__39_i800_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__39_i800_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__39_i800_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__39_i800_stall_in = 1'b0;
assign rnode_169to170_bb2__39_i800_0_NO_SHIFT_REG = rnode_169to170_bb2__39_i800_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__39_i800_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i800_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_or581_i788_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_valid_out_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_stall_in_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_or581_i788_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_or581_i788_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_or581_i788_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_or581_i788_0_stall_in_0_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_or581_i788_0_valid_out_0_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_or581_i788_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_or581_i788),
	.data_out(rnode_169to170_bb2_or581_i788_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_or581_i788_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_or581_i788_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_or581_i788_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_or581_i788_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_or581_i788_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or581_i788_stall_in = 1'b0;
assign rnode_169to170_bb2_or581_i788_0_stall_in_0_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i788_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2_or581_i788_0_NO_SHIFT_REG = rnode_169to170_bb2_or581_i788_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_or581_i788_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2_or581_i788_1_NO_SHIFT_REG = rnode_169to170_bb2_or581_i788_0_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and74_i794_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i794_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and74_i794_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i794_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and74_i794_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i794_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i794_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and74_i794_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and74_i794_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and74_i794_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and74_i794_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and74_i794_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and74_i794_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and74_i794),
	.data_out(rnode_169to170_bb2_and74_i794_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and74_i794_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and74_i794_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and74_i794_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and74_i794_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and74_i794_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and74_i794_stall_in = 1'b0;
assign rnode_169to170_bb2_and74_i794_0_NO_SHIFT_REG = rnode_169to170_bb2_and74_i794_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and74_i794_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and74_i794_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_cmp77_i333_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i333_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i333_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i333_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i333_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i333_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i333_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_cmp77_i333_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_cmp77_i333_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_cmp77_i333_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_cmp77_i333_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_cmp77_i333_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_cmp77_i333_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_cmp77_i333),
	.data_out(rnode_169to170_bb2_cmp77_i333_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_cmp77_i333_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_cmp77_i333_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2_cmp77_i333_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_cmp77_i333_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_cmp77_i333_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp77_i333_stall_in = 1'b0;
assign rnode_169to170_bb2_cmp77_i333_0_NO_SHIFT_REG = rnode_169to170_bb2_cmp77_i333_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_cmp77_i333_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i333_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__37_i322_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i322_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i322_1_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i322_2_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i322_3_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2__37_i322_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_valid_out_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_stall_in_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__37_i322_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__37_i322_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__37_i322_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__37_i322_0_stall_in_0_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__37_i322_0_valid_out_0_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__37_i322_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__37_i322),
	.data_out(rnode_169to170_bb2__37_i322_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__37_i322_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__37_i322_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2__37_i322_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__37_i322_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__37_i322_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__37_i322_stall_in = 1'b0;
assign rnode_169to170_bb2__37_i322_0_stall_in_0_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i322_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i322_0_NO_SHIFT_REG = rnode_169to170_bb2__37_i322_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i322_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i322_1_NO_SHIFT_REG = rnode_169to170_bb2__37_i322_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i322_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i322_2_NO_SHIFT_REG = rnode_169to170_bb2__37_i322_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__37_i322_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_169to170_bb2__37_i322_3_NO_SHIFT_REG = rnode_169to170_bb2__37_i322_0_reg_170_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2_and75_i328_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i328_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i328_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i328_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_169to170_bb2_and75_i328_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i328_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i328_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2_and75_i328_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2_and75_i328_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2_and75_i328_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2_and75_i328_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2_and75_i328_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2_and75_i328_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2_and75_i328),
	.data_out(rnode_169to170_bb2_and75_i328_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2_and75_i328_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2_and75_i328_0_reg_170_fifo.DATA_WIDTH = 32;
defparam rnode_169to170_bb2_and75_i328_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2_and75_i328_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2_and75_i328_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and75_i328_stall_in = 1'b0;
assign rnode_169to170_bb2_and75_i328_0_NO_SHIFT_REG = rnode_169to170_bb2_and75_i328_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2_and75_i328_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i328_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_169to170_bb2__39_i336_0_valid_out_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i336_0_stall_in_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i336_0_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i336_0_reg_170_inputs_ready_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i336_0_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i336_0_valid_out_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i336_0_stall_in_reg_170_NO_SHIFT_REG;
 logic rnode_169to170_bb2__39_i336_0_stall_out_reg_170_NO_SHIFT_REG;

acl_data_fifo rnode_169to170_bb2__39_i336_0_reg_170_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_169to170_bb2__39_i336_0_reg_170_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_169to170_bb2__39_i336_0_stall_in_reg_170_NO_SHIFT_REG),
	.valid_out(rnode_169to170_bb2__39_i336_0_valid_out_reg_170_NO_SHIFT_REG),
	.stall_out(rnode_169to170_bb2__39_i336_0_stall_out_reg_170_NO_SHIFT_REG),
	.data_in(local_bb2__39_i336),
	.data_out(rnode_169to170_bb2__39_i336_0_reg_170_NO_SHIFT_REG)
);

defparam rnode_169to170_bb2__39_i336_0_reg_170_fifo.DEPTH = 1;
defparam rnode_169to170_bb2__39_i336_0_reg_170_fifo.DATA_WIDTH = 1;
defparam rnode_169to170_bb2__39_i336_0_reg_170_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_169to170_bb2__39_i336_0_reg_170_fifo.IMPL = "shift_reg";

assign rnode_169to170_bb2__39_i336_0_reg_170_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__39_i336_stall_in = 1'b0;
assign rnode_169to170_bb2__39_i336_0_NO_SHIFT_REG = rnode_169to170_bb2__39_i336_0_reg_170_NO_SHIFT_REG;
assign rnode_169to170_bb2__39_i336_0_stall_in_reg_170_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i336_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u86_stall_local;
wire [31:0] local_bb2_var__u86;

assign local_bb2_var__u86[31:1] = 31'h0;
assign local_bb2_var__u86[0] = rnode_169to170_bb2_cmp68_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__40_i_stall_local;
wire local_bb2__40_i;

assign local_bb2__40_i = (rnode_169to170_bb2_cmp77_i_0_NO_SHIFT_REG | rnode_169to170_bb2__39_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i_stall_local;
wire local_bb2_reduction_2_i;

assign local_bb2_reduction_2_i = (rnode_169to170_bb2_reduction_0_i_0_NO_SHIFT_REG | rnode_169to170_bb2_or581_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cond111_i_stall_local;
wire [31:0] local_bb2_cond111_i;

assign local_bb2_cond111_i = (rnode_169to170_bb2_or581_i_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i_stall_local;
wire [31:0] local_bb2_shl_i;

assign local_bb2_shl_i = (rnode_169to170_bb2_and74_i_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp53_i1427_stall_local;
wire local_bb2_cmp53_i1427;

assign local_bb2_cmp53_i1427 = (rnode_169to170_bb2__37_i1426_0_NO_SHIFT_REG > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp68_i1431_stall_local;
wire local_bb2_cmp68_i1431;

assign local_bb2_cmp68_i1431 = (rnode_169to170_bb2__37_i1426_1_NO_SHIFT_REG < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i1433_stall_local;
wire [31:0] local_bb2_sub_i1433;

assign local_bb2_sub_i1433 = (rnode_169to170_bb2__37_i1426_2_NO_SHIFT_REG << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp71_not_i1448_stall_local;
wire local_bb2_cmp71_not_i1448;

assign local_bb2_cmp71_not_i1448 = (rnode_169to170_bb2__37_i1426_3_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__40_i1441_stall_local;
wire local_bb2__40_i1441;

assign local_bb2__40_i1441 = (rnode_169to170_bb2_cmp77_i1437_0_NO_SHIFT_REG | rnode_169to170_bb2__39_i1440_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp53_i879_stall_local;
wire local_bb2_cmp53_i879;

assign local_bb2_cmp53_i879 = (rnode_169to170_bb2__37_i878_0_NO_SHIFT_REG > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp68_i883_stall_local;
wire local_bb2_cmp68_i883;

assign local_bb2_cmp68_i883 = (rnode_169to170_bb2__37_i878_1_NO_SHIFT_REG < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i885_stall_local;
wire [31:0] local_bb2_sub_i885;

assign local_bb2_sub_i885 = (rnode_169to170_bb2__37_i878_2_NO_SHIFT_REG << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp71_not_i900_stall_local;
wire local_bb2_cmp71_not_i900;

assign local_bb2_cmp71_not_i900 = (rnode_169to170_bb2__37_i878_3_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__40_i893_stall_local;
wire local_bb2__40_i893;

assign local_bb2__40_i893 = (rnode_169to170_bb2_cmp77_i889_0_NO_SHIFT_REG | rnode_169to170_bb2__39_i892_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp53_i415_stall_local;
wire local_bb2_cmp53_i415;

assign local_bb2_cmp53_i415 = (rnode_169to170_bb2__37_i414_0_NO_SHIFT_REG > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp68_i419_stall_local;
wire local_bb2_cmp68_i419;

assign local_bb2_cmp68_i419 = (rnode_169to170_bb2__37_i414_1_NO_SHIFT_REG < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i421_stall_local;
wire [31:0] local_bb2_sub_i421;

assign local_bb2_sub_i421 = (rnode_169to170_bb2__37_i414_2_NO_SHIFT_REG << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp71_not_i436_stall_local;
wire local_bb2_cmp71_not_i436;

assign local_bb2_cmp71_not_i436 = (rnode_169to170_bb2__37_i414_3_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__40_i429_stall_local;
wire local_bb2__40_i429;

assign local_bb2__40_i429 = (rnode_169to170_bb2_cmp77_i425_0_NO_SHIFT_REG | rnode_169to170_bb2__39_i428_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u87_stall_local;
wire [31:0] local_bb2_var__u87;

assign local_bb2_var__u87[31:1] = 31'h0;
assign local_bb2_var__u87[0] = rnode_169to170_bb2_cmp68_i1888_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__40_i1898_stall_local;
wire local_bb2__40_i1898;

assign local_bb2__40_i1898 = (rnode_169to170_bb2_cmp77_i1894_0_NO_SHIFT_REG | rnode_169to170_bb2__39_i1897_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i1887_stall_local;
wire local_bb2_reduction_2_i1887;

assign local_bb2_reduction_2_i1887 = (rnode_169to170_bb2_reduction_0_i1886_0_NO_SHIFT_REG | rnode_169to170_bb2_or581_i1885_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cond111_i1913_stall_local;
wire [31:0] local_bb2_cond111_i1913;

assign local_bb2_cond111_i1913 = (rnode_169to170_bb2_or581_i1885_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i1892_stall_local;
wire [31:0] local_bb2_shl_i1892;

assign local_bb2_shl_i1892 = (rnode_169to170_bb2_and74_i1891_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp53_i1335_stall_local;
wire local_bb2_cmp53_i1335;

assign local_bb2_cmp53_i1335 = (rnode_169to170_bb2__37_i1334_0_NO_SHIFT_REG > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp68_i1339_stall_local;
wire local_bb2_cmp68_i1339;

assign local_bb2_cmp68_i1339 = (rnode_169to170_bb2__37_i1334_1_NO_SHIFT_REG < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i1341_stall_local;
wire [31:0] local_bb2_sub_i1341;

assign local_bb2_sub_i1341 = (rnode_169to170_bb2__37_i1334_2_NO_SHIFT_REG << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp71_not_i1356_stall_local;
wire local_bb2_cmp71_not_i1356;

assign local_bb2_cmp71_not_i1356 = (rnode_169to170_bb2__37_i1334_3_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__40_i1349_stall_local;
wire local_bb2__40_i1349;

assign local_bb2__40_i1349 = (rnode_169to170_bb2_cmp77_i1345_0_NO_SHIFT_REG | rnode_169to170_bb2__39_i1348_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u88_stall_local;
wire [31:0] local_bb2_var__u88;

assign local_bb2_var__u88[31:1] = 31'h0;
assign local_bb2_var__u88[0] = rnode_169to170_bb2_cmp68_i791_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__40_i801_stall_local;
wire local_bb2__40_i801;

assign local_bb2__40_i801 = (rnode_169to170_bb2_cmp77_i797_0_NO_SHIFT_REG | rnode_169to170_bb2__39_i800_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i790_stall_local;
wire local_bb2_reduction_2_i790;

assign local_bb2_reduction_2_i790 = (rnode_169to170_bb2_reduction_0_i789_0_NO_SHIFT_REG | rnode_169to170_bb2_or581_i788_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cond111_i816_stall_local;
wire [31:0] local_bb2_cond111_i816;

assign local_bb2_cond111_i816 = (rnode_169to170_bb2_or581_i788_1_NO_SHIFT_REG ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i795_stall_local;
wire [31:0] local_bb2_shl_i795;

assign local_bb2_shl_i795 = (rnode_169to170_bb2_and74_i794_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp53_i323_stall_local;
wire local_bb2_cmp53_i323;

assign local_bb2_cmp53_i323 = (rnode_169to170_bb2__37_i322_0_NO_SHIFT_REG > 32'h17D);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp68_i327_stall_local;
wire local_bb2_cmp68_i327;

assign local_bb2_cmp68_i327 = (rnode_169to170_bb2__37_i322_1_NO_SHIFT_REG < 32'h80);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i329_stall_local;
wire [31:0] local_bb2_sub_i329;

assign local_bb2_sub_i329 = (rnode_169to170_bb2__37_i322_2_NO_SHIFT_REG << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp71_not_i344_stall_local;
wire local_bb2_cmp71_not_i344;

assign local_bb2_cmp71_not_i344 = (rnode_169to170_bb2__37_i322_3_NO_SHIFT_REG != 32'h7F);

// This section implements an unregistered operation.
// 
wire local_bb2__40_i337_stall_local;
wire local_bb2__40_i337;

assign local_bb2__40_i337 = (rnode_169to170_bb2_cmp77_i333_0_NO_SHIFT_REG | rnode_169to170_bb2__39_i336_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cond_i_stall_local;
wire [31:0] local_bb2_cond_i;

assign local_bb2_cond_i[31:1] = 31'h0;
assign local_bb2_cond_i[0] = local_bb2__40_i;

// This section implements an unregistered operation.
// 
wire local_bb2_conv101_i_stall_local;
wire [31:0] local_bb2_conv101_i;

assign local_bb2_conv101_i[31:1] = 31'h0;
assign local_bb2_conv101_i[0] = local_bb2_reduction_2_i;

// This section implements an unregistered operation.
// 
wire local_bb2_or76_i_stall_local;
wire [31:0] local_bb2_or76_i;

assign local_bb2_or76_i = (local_bb2_shl_i | rnode_169to170_bb2_and75_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_or581_i1428_stall_local;
wire local_bb2_or581_i1428;

assign local_bb2_or581_i1428 = (rnode_169to170_bb2_var__u48_0_NO_SHIFT_REG | local_bb2_cmp53_i1427);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u89_stall_local;
wire [31:0] local_bb2_var__u89;

assign local_bb2_var__u89[31:1] = 31'h0;
assign local_bb2_var__u89[0] = local_bb2_cmp68_i1431;

// This section implements an unregistered operation.
// 
wire local_bb2_and74_i1434_stall_local;
wire [31:0] local_bb2_and74_i1434;

assign local_bb2_and74_i1434 = (local_bb2_sub_i1433 + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cond_i1442_stall_local;
wire [31:0] local_bb2_cond_i1442;

assign local_bb2_cond_i1442[31:1] = 31'h0;
assign local_bb2_cond_i1442[0] = local_bb2__40_i1441;

// This section implements an unregistered operation.
// 
wire local_bb2_or581_i880_stall_local;
wire local_bb2_or581_i880;

assign local_bb2_or581_i880 = (rnode_169to170_bb2_var__u50_0_NO_SHIFT_REG | local_bb2_cmp53_i879);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u90_stall_local;
wire [31:0] local_bb2_var__u90;

assign local_bb2_var__u90[31:1] = 31'h0;
assign local_bb2_var__u90[0] = local_bb2_cmp68_i883;

// This section implements an unregistered operation.
// 
wire local_bb2_and74_i886_stall_local;
wire [31:0] local_bb2_and74_i886;

assign local_bb2_and74_i886 = (local_bb2_sub_i885 + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cond_i894_stall_local;
wire [31:0] local_bb2_cond_i894;

assign local_bb2_cond_i894[31:1] = 31'h0;
assign local_bb2_cond_i894[0] = local_bb2__40_i893;

// This section implements an unregistered operation.
// 
wire local_bb2_or581_i416_stall_local;
wire local_bb2_or581_i416;

assign local_bb2_or581_i416 = (rnode_169to170_bb2_var__u52_0_NO_SHIFT_REG | local_bb2_cmp53_i415);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u91_stall_local;
wire [31:0] local_bb2_var__u91;

assign local_bb2_var__u91[31:1] = 31'h0;
assign local_bb2_var__u91[0] = local_bb2_cmp68_i419;

// This section implements an unregistered operation.
// 
wire local_bb2_and74_i422_stall_local;
wire [31:0] local_bb2_and74_i422;

assign local_bb2_and74_i422 = (local_bb2_sub_i421 + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cond_i430_stall_local;
wire [31:0] local_bb2_cond_i430;

assign local_bb2_cond_i430[31:1] = 31'h0;
assign local_bb2_cond_i430[0] = local_bb2__40_i429;

// This section implements an unregistered operation.
// 
wire local_bb2_cond_i1899_stall_local;
wire [31:0] local_bb2_cond_i1899;

assign local_bb2_cond_i1899[31:1] = 31'h0;
assign local_bb2_cond_i1899[0] = local_bb2__40_i1898;

// This section implements an unregistered operation.
// 
wire local_bb2_conv101_i1908_stall_local;
wire [31:0] local_bb2_conv101_i1908;

assign local_bb2_conv101_i1908[31:1] = 31'h0;
assign local_bb2_conv101_i1908[0] = local_bb2_reduction_2_i1887;

// This section implements an unregistered operation.
// 
wire local_bb2_or76_i1893_stall_local;
wire [31:0] local_bb2_or76_i1893;

assign local_bb2_or76_i1893 = (local_bb2_shl_i1892 | rnode_169to170_bb2_and75_i1889_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_or581_i1336_stall_local;
wire local_bb2_or581_i1336;

assign local_bb2_or581_i1336 = (rnode_169to170_bb2_var__u56_0_NO_SHIFT_REG | local_bb2_cmp53_i1335);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u92_stall_local;
wire [31:0] local_bb2_var__u92;

assign local_bb2_var__u92[31:1] = 31'h0;
assign local_bb2_var__u92[0] = local_bb2_cmp68_i1339;

// This section implements an unregistered operation.
// 
wire local_bb2_and74_i1342_stall_local;
wire [31:0] local_bb2_and74_i1342;

assign local_bb2_and74_i1342 = (local_bb2_sub_i1341 + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cond_i1350_stall_local;
wire [31:0] local_bb2_cond_i1350;

assign local_bb2_cond_i1350[31:1] = 31'h0;
assign local_bb2_cond_i1350[0] = local_bb2__40_i1349;

// This section implements an unregistered operation.
// 
wire local_bb2_cond_i802_stall_local;
wire [31:0] local_bb2_cond_i802;

assign local_bb2_cond_i802[31:1] = 31'h0;
assign local_bb2_cond_i802[0] = local_bb2__40_i801;

// This section implements an unregistered operation.
// 
wire local_bb2_conv101_i811_stall_local;
wire [31:0] local_bb2_conv101_i811;

assign local_bb2_conv101_i811[31:1] = 31'h0;
assign local_bb2_conv101_i811[0] = local_bb2_reduction_2_i790;

// This section implements an unregistered operation.
// 
wire local_bb2_or76_i796_stall_local;
wire [31:0] local_bb2_or76_i796;

assign local_bb2_or76_i796 = (local_bb2_shl_i795 | rnode_169to170_bb2_and75_i792_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_or581_i324_stall_local;
wire local_bb2_or581_i324;

assign local_bb2_or581_i324 = (rnode_169to170_bb2_var__u60_0_NO_SHIFT_REG | local_bb2_cmp53_i323);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u93_stall_local;
wire [31:0] local_bb2_var__u93;

assign local_bb2_var__u93[31:1] = 31'h0;
assign local_bb2_var__u93[0] = local_bb2_cmp68_i327;

// This section implements an unregistered operation.
// 
wire local_bb2_and74_i330_stall_local;
wire [31:0] local_bb2_and74_i330;

assign local_bb2_and74_i330 = (local_bb2_sub_i329 + 32'h40800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cond_i338_stall_local;
wire [31:0] local_bb2_cond_i338;

assign local_bb2_cond_i338[31:1] = 31'h0;
assign local_bb2_cond_i338[0] = local_bb2__40_i337;

// This section implements an unregistered operation.
// 
wire local_bb2_add87_i_stall_local;
wire [31:0] local_bb2_add87_i;

assign local_bb2_add87_i = (local_bb2_cond_i + local_bb2_or76_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i1430_stall_local;
wire local_bb2_reduction_2_i1430;

assign local_bb2_reduction_2_i1430 = (rnode_169to170_bb2_reduction_0_i1429_0_NO_SHIFT_REG | local_bb2_or581_i1428);

// This section implements an unregistered operation.
// 
wire local_bb2_cond111_i1456_stall_local;
wire [31:0] local_bb2_cond111_i1456;

assign local_bb2_cond111_i1456 = (local_bb2_or581_i1428 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i1435_stall_local;
wire [31:0] local_bb2_shl_i1435;

assign local_bb2_shl_i1435 = (local_bb2_and74_i1434 & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i882_stall_local;
wire local_bb2_reduction_2_i882;

assign local_bb2_reduction_2_i882 = (rnode_169to170_bb2_reduction_0_i881_0_NO_SHIFT_REG | local_bb2_or581_i880);

// This section implements an unregistered operation.
// 
wire local_bb2_cond111_i908_stall_local;
wire [31:0] local_bb2_cond111_i908;

assign local_bb2_cond111_i908 = (local_bb2_or581_i880 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i887_stall_local;
wire [31:0] local_bb2_shl_i887;

assign local_bb2_shl_i887 = (local_bb2_and74_i886 & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i418_stall_local;
wire local_bb2_reduction_2_i418;

assign local_bb2_reduction_2_i418 = (rnode_169to170_bb2_reduction_0_i417_0_NO_SHIFT_REG | local_bb2_or581_i416);

// This section implements an unregistered operation.
// 
wire local_bb2_cond111_i444_stall_local;
wire [31:0] local_bb2_cond111_i444;

assign local_bb2_cond111_i444 = (local_bb2_or581_i416 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i423_stall_local;
wire [31:0] local_bb2_shl_i423;

assign local_bb2_shl_i423 = (local_bb2_and74_i422 & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_add87_i1900_stall_local;
wire [31:0] local_bb2_add87_i1900;

assign local_bb2_add87_i1900 = (local_bb2_cond_i1899 + local_bb2_or76_i1893);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i1338_stall_local;
wire local_bb2_reduction_2_i1338;

assign local_bb2_reduction_2_i1338 = (rnode_169to170_bb2_reduction_0_i1337_0_NO_SHIFT_REG | local_bb2_or581_i1336);

// This section implements an unregistered operation.
// 
wire local_bb2_cond111_i1364_stall_local;
wire [31:0] local_bb2_cond111_i1364;

assign local_bb2_cond111_i1364 = (local_bb2_or581_i1336 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i1343_stall_local;
wire [31:0] local_bb2_shl_i1343;

assign local_bb2_shl_i1343 = (local_bb2_and74_i1342 & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_add87_i803_stall_local;
wire [31:0] local_bb2_add87_i803;

assign local_bb2_add87_i803 = (local_bb2_cond_i802 + local_bb2_or76_i796);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i326_stall_local;
wire local_bb2_reduction_2_i326;

assign local_bb2_reduction_2_i326 = (rnode_169to170_bb2_reduction_0_i325_0_NO_SHIFT_REG | local_bb2_or581_i324);

// This section implements an unregistered operation.
// 
wire local_bb2_cond111_i352_stall_local;
wire [31:0] local_bb2_cond111_i352;

assign local_bb2_cond111_i352 = (local_bb2_or581_i324 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i331_stall_local;
wire [31:0] local_bb2_shl_i331;

assign local_bb2_shl_i331 = (local_bb2_and74_i330 & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i_stall_local;
wire [31:0] local_bb2_and88_i;

assign local_bb2_and88_i = (local_bb2_add87_i & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i_stall_local;
wire [31:0] local_bb2_and90_i;

assign local_bb2_and90_i = (local_bb2_add87_i & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_conv101_i1451_stall_local;
wire [31:0] local_bb2_conv101_i1451;

assign local_bb2_conv101_i1451[31:1] = 31'h0;
assign local_bb2_conv101_i1451[0] = local_bb2_reduction_2_i1430;

// This section implements an unregistered operation.
// 
wire local_bb2_or76_i1436_stall_local;
wire [31:0] local_bb2_or76_i1436;

assign local_bb2_or76_i1436 = (local_bb2_shl_i1435 | rnode_169to170_bb2_and75_i1432_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_conv101_i903_stall_local;
wire [31:0] local_bb2_conv101_i903;

assign local_bb2_conv101_i903[31:1] = 31'h0;
assign local_bb2_conv101_i903[0] = local_bb2_reduction_2_i882;

// This section implements an unregistered operation.
// 
wire local_bb2_or76_i888_stall_local;
wire [31:0] local_bb2_or76_i888;

assign local_bb2_or76_i888 = (local_bb2_shl_i887 | rnode_169to170_bb2_and75_i884_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_conv101_i439_stall_local;
wire [31:0] local_bb2_conv101_i439;

assign local_bb2_conv101_i439[31:1] = 31'h0;
assign local_bb2_conv101_i439[0] = local_bb2_reduction_2_i418;

// This section implements an unregistered operation.
// 
wire local_bb2_or76_i424_stall_local;
wire [31:0] local_bb2_or76_i424;

assign local_bb2_or76_i424 = (local_bb2_shl_i423 | rnode_169to170_bb2_and75_i420_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i1901_stall_local;
wire [31:0] local_bb2_and88_i1901;

assign local_bb2_and88_i1901 = (local_bb2_add87_i1900 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i1903_stall_local;
wire [31:0] local_bb2_and90_i1903;

assign local_bb2_and90_i1903 = (local_bb2_add87_i1900 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_conv101_i1359_stall_local;
wire [31:0] local_bb2_conv101_i1359;

assign local_bb2_conv101_i1359[31:1] = 31'h0;
assign local_bb2_conv101_i1359[0] = local_bb2_reduction_2_i1338;

// This section implements an unregistered operation.
// 
wire local_bb2_or76_i1344_stall_local;
wire [31:0] local_bb2_or76_i1344;

assign local_bb2_or76_i1344 = (local_bb2_shl_i1343 | rnode_169to170_bb2_and75_i1340_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i804_stall_local;
wire [31:0] local_bb2_and88_i804;

assign local_bb2_and88_i804 = (local_bb2_add87_i803 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i806_stall_local;
wire [31:0] local_bb2_and90_i806;

assign local_bb2_and90_i806 = (local_bb2_add87_i803 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_conv101_i347_stall_local;
wire [31:0] local_bb2_conv101_i347;

assign local_bb2_conv101_i347[31:1] = 31'h0;
assign local_bb2_conv101_i347[0] = local_bb2_reduction_2_i326;

// This section implements an unregistered operation.
// 
wire local_bb2_or76_i332_stall_local;
wire [31:0] local_bb2_or76_i332;

assign local_bb2_or76_i332 = (local_bb2_shl_i331 | rnode_169to170_bb2_and75_i328_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_or89_i_stall_local;
wire [31:0] local_bb2_or89_i;

assign local_bb2_or89_i = (local_bb2_and88_i | local_bb2_and4_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i_stall_local;
wire local_bb2_cmp91_i;

assign local_bb2_cmp91_i = (local_bb2_and90_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_add87_i1443_stall_local;
wire [31:0] local_bb2_add87_i1443;

assign local_bb2_add87_i1443 = (local_bb2_cond_i1442 + local_bb2_or76_i1436);

// This section implements an unregistered operation.
// 
wire local_bb2_add87_i895_stall_local;
wire [31:0] local_bb2_add87_i895;

assign local_bb2_add87_i895 = (local_bb2_cond_i894 + local_bb2_or76_i888);

// This section implements an unregistered operation.
// 
wire local_bb2_add87_i431_stall_local;
wire [31:0] local_bb2_add87_i431;

assign local_bb2_add87_i431 = (local_bb2_cond_i430 + local_bb2_or76_i424);

// This section implements an unregistered operation.
// 
wire local_bb2_or89_i1902_stall_local;
wire [31:0] local_bb2_or89_i1902;

assign local_bb2_or89_i1902 = (local_bb2_and88_i1901 | local_bb2_and4_i1828);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i1904_stall_local;
wire local_bb2_cmp91_i1904;

assign local_bb2_cmp91_i1904 = (local_bb2_and90_i1903 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_add87_i1351_stall_local;
wire [31:0] local_bb2_add87_i1351;

assign local_bb2_add87_i1351 = (local_bb2_cond_i1350 + local_bb2_or76_i1344);

// This section implements an unregistered operation.
// 
wire local_bb2_or89_i805_stall_local;
wire [31:0] local_bb2_or89_i805;

assign local_bb2_or89_i805 = (local_bb2_and88_i804 | local_bb2_and4_i731);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i807_stall_local;
wire local_bb2_cmp91_i807;

assign local_bb2_cmp91_i807 = (local_bb2_and90_i806 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_add87_i339_stall_local;
wire [31:0] local_bb2_add87_i339;

assign local_bb2_add87_i339 = (local_bb2_cond_i338 + local_bb2_or76_i332);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge14_i_stall_local;
wire local_bb2_brmerge14_i;

assign local_bb2_brmerge14_i = (local_bb2_cmp91_i | rnode_169to170_bb2_cmp71_not_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i1444_stall_local;
wire [31:0] local_bb2_and88_i1444;

assign local_bb2_and88_i1444 = (local_bb2_add87_i1443 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i1446_stall_local;
wire [31:0] local_bb2_and90_i1446;

assign local_bb2_and90_i1446 = (local_bb2_add87_i1443 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i896_stall_local;
wire [31:0] local_bb2_and88_i896;

assign local_bb2_and88_i896 = (local_bb2_add87_i895 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i898_stall_local;
wire [31:0] local_bb2_and90_i898;

assign local_bb2_and90_i898 = (local_bb2_add87_i895 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i432_stall_local;
wire [31:0] local_bb2_and88_i432;

assign local_bb2_and88_i432 = (local_bb2_add87_i431 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i434_stall_local;
wire [31:0] local_bb2_and90_i434;

assign local_bb2_and90_i434 = (local_bb2_add87_i431 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge14_i1906_stall_local;
wire local_bb2_brmerge14_i1906;

assign local_bb2_brmerge14_i1906 = (local_bb2_cmp91_i1904 | rnode_169to170_bb2_cmp71_not_i1905_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i1352_stall_local;
wire [31:0] local_bb2_and88_i1352;

assign local_bb2_and88_i1352 = (local_bb2_add87_i1351 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i1354_stall_local;
wire [31:0] local_bb2_and90_i1354;

assign local_bb2_and90_i1354 = (local_bb2_add87_i1351 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge14_i809_stall_local;
wire local_bb2_brmerge14_i809;

assign local_bb2_brmerge14_i809 = (local_bb2_cmp91_i807 | rnode_169to170_bb2_cmp71_not_i808_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i340_stall_local;
wire [31:0] local_bb2_and88_i340;

assign local_bb2_and88_i340 = (local_bb2_add87_i339 & 32'h7FFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i342_stall_local;
wire [31:0] local_bb2_and90_i342;

assign local_bb2_and90_i342 = (local_bb2_add87_i339 & 32'h800000);

// This section implements an unregistered operation.
// 
wire local_bb2_conv99_i_stall_local;
wire [31:0] local_bb2_conv99_i;

assign local_bb2_conv99_i = (local_bb2_brmerge14_i ? local_bb2_var__u86 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or89_i1445_stall_local;
wire [31:0] local_bb2_or89_i1445;

assign local_bb2_or89_i1445 = (local_bb2_and88_i1444 | local_bb2_and4_i1371);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i1447_stall_local;
wire local_bb2_cmp91_i1447;

assign local_bb2_cmp91_i1447 = (local_bb2_and90_i1446 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or89_i897_stall_local;
wire [31:0] local_bb2_or89_i897;

assign local_bb2_or89_i897 = (local_bb2_and88_i896 | local_bb2_and4_i823);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i899_stall_local;
wire local_bb2_cmp91_i899;

assign local_bb2_cmp91_i899 = (local_bb2_and90_i898 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or89_i433_stall_local;
wire [31:0] local_bb2_or89_i433;

assign local_bb2_or89_i433 = (local_bb2_and88_i432 | local_bb2_and4_i359);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i435_stall_local;
wire local_bb2_cmp91_i435;

assign local_bb2_cmp91_i435 = (local_bb2_and90_i434 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_conv99_i1907_stall_local;
wire [31:0] local_bb2_conv99_i1907;

assign local_bb2_conv99_i1907 = (local_bb2_brmerge14_i1906 ? local_bb2_var__u87 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or89_i1353_stall_local;
wire [31:0] local_bb2_or89_i1353;

assign local_bb2_or89_i1353 = (local_bb2_and88_i1352 | local_bb2_and4_i1279);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i1355_stall_local;
wire local_bb2_cmp91_i1355;

assign local_bb2_cmp91_i1355 = (local_bb2_and90_i1354 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_conv99_i810_stall_local;
wire [31:0] local_bb2_conv99_i810;

assign local_bb2_conv99_i810 = (local_bb2_brmerge14_i809 ? local_bb2_var__u88 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or89_i341_stall_local;
wire [31:0] local_bb2_or89_i341;

assign local_bb2_or89_i341 = (local_bb2_and88_i340 | local_bb2_and4_i267);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i343_stall_local;
wire local_bb2_cmp91_i343;

assign local_bb2_cmp91_i343 = (local_bb2_and90_i342 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or102_i_stall_local;
wire [31:0] local_bb2_or102_i;

assign local_bb2_or102_i = (local_bb2_conv99_i | local_bb2_conv101_i);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge14_i1449_stall_local;
wire local_bb2_brmerge14_i1449;

assign local_bb2_brmerge14_i1449 = (local_bb2_cmp91_i1447 | local_bb2_cmp71_not_i1448);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge14_i901_stall_local;
wire local_bb2_brmerge14_i901;

assign local_bb2_brmerge14_i901 = (local_bb2_cmp91_i899 | local_bb2_cmp71_not_i900);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge14_i437_stall_local;
wire local_bb2_brmerge14_i437;

assign local_bb2_brmerge14_i437 = (local_bb2_cmp91_i435 | local_bb2_cmp71_not_i436);

// This section implements an unregistered operation.
// 
wire local_bb2_or102_i1909_stall_local;
wire [31:0] local_bb2_or102_i1909;

assign local_bb2_or102_i1909 = (local_bb2_conv99_i1907 | local_bb2_conv101_i1908);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge14_i1357_stall_local;
wire local_bb2_brmerge14_i1357;

assign local_bb2_brmerge14_i1357 = (local_bb2_cmp91_i1355 | local_bb2_cmp71_not_i1356);

// This section implements an unregistered operation.
// 
wire local_bb2_or102_i812_stall_local;
wire [31:0] local_bb2_or102_i812;

assign local_bb2_or102_i812 = (local_bb2_conv99_i810 | local_bb2_conv101_i811);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge14_i345_stall_local;
wire local_bb2_brmerge14_i345;

assign local_bb2_brmerge14_i345 = (local_bb2_cmp91_i343 | local_bb2_cmp71_not_i344);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool103_i_stall_local;
wire local_bb2_tobool103_i;

assign local_bb2_tobool103_i = (local_bb2_or102_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_conv99_i1450_stall_local;
wire [31:0] local_bb2_conv99_i1450;

assign local_bb2_conv99_i1450 = (local_bb2_brmerge14_i1449 ? local_bb2_var__u89 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_conv99_i902_stall_local;
wire [31:0] local_bb2_conv99_i902;

assign local_bb2_conv99_i902 = (local_bb2_brmerge14_i901 ? local_bb2_var__u90 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_conv99_i438_stall_local;
wire [31:0] local_bb2_conv99_i438;

assign local_bb2_conv99_i438 = (local_bb2_brmerge14_i437 ? local_bb2_var__u91 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool103_i1910_stall_local;
wire local_bb2_tobool103_i1910;

assign local_bb2_tobool103_i1910 = (local_bb2_or102_i1909 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_conv99_i1358_stall_local;
wire [31:0] local_bb2_conv99_i1358;

assign local_bb2_conv99_i1358 = (local_bb2_brmerge14_i1357 ? local_bb2_var__u92 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool103_i813_stall_local;
wire local_bb2_tobool103_i813;

assign local_bb2_tobool103_i813 = (local_bb2_or102_i812 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_conv99_i346_stall_local;
wire [31:0] local_bb2_conv99_i346;

assign local_bb2_conv99_i346 = (local_bb2_brmerge14_i345 ? local_bb2_var__u93 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cond107_i_stall_local;
wire [31:0] local_bb2_cond107_i;

assign local_bb2_cond107_i = (local_bb2_tobool103_i ? local_bb2_and4_i : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or102_i1452_stall_local;
wire [31:0] local_bb2_or102_i1452;

assign local_bb2_or102_i1452 = (local_bb2_conv99_i1450 | local_bb2_conv101_i1451);

// This section implements an unregistered operation.
// 
wire local_bb2_or102_i904_stall_local;
wire [31:0] local_bb2_or102_i904;

assign local_bb2_or102_i904 = (local_bb2_conv99_i902 | local_bb2_conv101_i903);

// This section implements an unregistered operation.
// 
wire local_bb2_or102_i440_stall_local;
wire [31:0] local_bb2_or102_i440;

assign local_bb2_or102_i440 = (local_bb2_conv99_i438 | local_bb2_conv101_i439);

// This section implements an unregistered operation.
// 
wire local_bb2_cond107_i1911_stall_local;
wire [31:0] local_bb2_cond107_i1911;

assign local_bb2_cond107_i1911 = (local_bb2_tobool103_i1910 ? local_bb2_and4_i1828 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or102_i1360_stall_local;
wire [31:0] local_bb2_or102_i1360;

assign local_bb2_or102_i1360 = (local_bb2_conv99_i1358 | local_bb2_conv101_i1359);

// This section implements an unregistered operation.
// 
wire local_bb2_cond107_i814_stall_local;
wire [31:0] local_bb2_cond107_i814;

assign local_bb2_cond107_i814 = (local_bb2_tobool103_i813 ? local_bb2_and4_i731 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or102_i348_stall_local;
wire [31:0] local_bb2_or102_i348;

assign local_bb2_or102_i348 = (local_bb2_conv99_i346 | local_bb2_conv101_i347);

// This section implements an unregistered operation.
// 
wire local_bb2_and108_i_stall_local;
wire [31:0] local_bb2_and108_i;

assign local_bb2_and108_i = (local_bb2_cond107_i & local_bb2_or89_i);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool103_i1453_stall_local;
wire local_bb2_tobool103_i1453;

assign local_bb2_tobool103_i1453 = (local_bb2_or102_i1452 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool103_i905_stall_local;
wire local_bb2_tobool103_i905;

assign local_bb2_tobool103_i905 = (local_bb2_or102_i904 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool103_i441_stall_local;
wire local_bb2_tobool103_i441;

assign local_bb2_tobool103_i441 = (local_bb2_or102_i440 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_and108_i1912_stall_local;
wire [31:0] local_bb2_and108_i1912;

assign local_bb2_and108_i1912 = (local_bb2_cond107_i1911 & local_bb2_or89_i1902);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool103_i1361_stall_local;
wire local_bb2_tobool103_i1361;

assign local_bb2_tobool103_i1361 = (local_bb2_or102_i1360 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_and108_i815_stall_local;
wire [31:0] local_bb2_and108_i815;

assign local_bb2_and108_i815 = (local_bb2_cond107_i814 & local_bb2_or89_i805);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool103_i349_stall_local;
wire local_bb2_tobool103_i349;

assign local_bb2_tobool103_i349 = (local_bb2_or102_i348 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i_stall_local;
wire [31:0] local_bb2_or112_i;

assign local_bb2_or112_i = (local_bb2_and108_i | local_bb2_cond111_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cond107_i1454_stall_local;
wire [31:0] local_bb2_cond107_i1454;

assign local_bb2_cond107_i1454 = (local_bb2_tobool103_i1453 ? local_bb2_and4_i1371 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond107_i906_stall_local;
wire [31:0] local_bb2_cond107_i906;

assign local_bb2_cond107_i906 = (local_bb2_tobool103_i905 ? local_bb2_and4_i823 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond107_i442_stall_local;
wire [31:0] local_bb2_cond107_i442;

assign local_bb2_cond107_i442 = (local_bb2_tobool103_i441 ? local_bb2_and4_i359 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i1914_stall_local;
wire [31:0] local_bb2_or112_i1914;

assign local_bb2_or112_i1914 = (local_bb2_and108_i1912 | local_bb2_cond111_i1913);

// This section implements an unregistered operation.
// 
wire local_bb2_cond107_i1362_stall_local;
wire [31:0] local_bb2_cond107_i1362;

assign local_bb2_cond107_i1362 = (local_bb2_tobool103_i1361 ? local_bb2_and4_i1279 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i817_stall_local;
wire [31:0] local_bb2_or112_i817;

assign local_bb2_or112_i817 = (local_bb2_and108_i815 | local_bb2_cond111_i816);

// This section implements an unregistered operation.
// 
wire local_bb2_cond107_i350_stall_local;
wire [31:0] local_bb2_cond107_i350;

assign local_bb2_cond107_i350 = (local_bb2_tobool103_i349 ? local_bb2_and4_i267 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u94_valid_out;
wire local_bb2_var__u94_stall_in;
wire local_bb2_var__u94_inputs_ready;
wire local_bb2_var__u94_stall_local;
wire [31:0] local_bb2_var__u94;

assign local_bb2_var__u94_inputs_ready = (rnode_169to170_bb2_xor_i_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__29_i_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_or581_i_0_valid_out_1_NO_SHIFT_REG & rnode_169to170_bb2_or581_i_0_valid_out_0_NO_SHIFT_REG & rnode_169to170_bb2_reduction_0_i_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp68_i_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp71_not_i_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp77_i_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__39_i_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and75_i_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and74_i_0_valid_out_NO_SHIFT_REG);
assign local_bb2_var__u94 = (rnode_169to170_bb2__29_i_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb2_or112_i);
assign local_bb2_var__u94_valid_out = 1'b1;
assign rnode_169to170_bb2_xor_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp68_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and74_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and108_i1455_stall_local;
wire [31:0] local_bb2_and108_i1455;

assign local_bb2_and108_i1455 = (local_bb2_cond107_i1454 & local_bb2_or89_i1445);

// This section implements an unregistered operation.
// 
wire local_bb2_and108_i907_stall_local;
wire [31:0] local_bb2_and108_i907;

assign local_bb2_and108_i907 = (local_bb2_cond107_i906 & local_bb2_or89_i897);

// This section implements an unregistered operation.
// 
wire local_bb2_and108_i443_stall_local;
wire [31:0] local_bb2_and108_i443;

assign local_bb2_and108_i443 = (local_bb2_cond107_i442 & local_bb2_or89_i433);

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i1914_op_stall_local;
wire [31:0] local_bb2_or112_i1914_op;

assign local_bb2_or112_i1914_op = (local_bb2_or112_i1914 ^ 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and108_i1363_stall_local;
wire [31:0] local_bb2_and108_i1363;

assign local_bb2_and108_i1363 = (local_bb2_cond107_i1362 & local_bb2_or89_i1353);

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i817_op_stall_local;
wire [31:0] local_bb2_or112_i817_op;

assign local_bb2_or112_i817_op = (local_bb2_or112_i817 ^ 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and108_i351_stall_local;
wire [31:0] local_bb2_and108_i351;

assign local_bb2_and108_i351 = (local_bb2_cond107_i350 & local_bb2_or89_i341);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb2_var__u94_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u94_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u94_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u94_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u94_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u94_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u94_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb2_var__u94_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb2_var__u94_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb2_var__u94_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb2_var__u94_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb2_var__u94_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb2_var__u94),
	.data_out(rnode_170to171_bb2_var__u94_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb2_var__u94_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_bb2_var__u94_0_reg_171_fifo.DATA_WIDTH = 32;
defparam rnode_170to171_bb2_var__u94_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_bb2_var__u94_0_reg_171_fifo.IMPL = "shift_reg";

assign rnode_170to171_bb2_var__u94_0_reg_171_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u94_stall_in = 1'b0;
assign rnode_170to171_bb2_var__u94_0_stall_in_0_reg_171_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u94_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u94_0_NO_SHIFT_REG = rnode_170to171_bb2_var__u94_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u94_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u94_1_NO_SHIFT_REG = rnode_170to171_bb2_var__u94_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u94_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u94_2_NO_SHIFT_REG = rnode_170to171_bb2_var__u94_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u94_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u94_3_NO_SHIFT_REG = rnode_170to171_bb2_var__u94_0_reg_171_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i1457_stall_local;
wire [31:0] local_bb2_or112_i1457;

assign local_bb2_or112_i1457 = (local_bb2_and108_i1455 | local_bb2_cond111_i1456);

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i909_stall_local;
wire [31:0] local_bb2_or112_i909;

assign local_bb2_or112_i909 = (local_bb2_and108_i907 | local_bb2_cond111_i908);

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i445_stall_local;
wire [31:0] local_bb2_or112_i445;

assign local_bb2_or112_i445 = (local_bb2_and108_i443 | local_bb2_cond111_i444);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i1640_valid_out;
wire local_bb2_xor_i1640_stall_in;
wire local_bb2_xor_i1640_inputs_ready;
wire local_bb2_xor_i1640_stall_local;
wire [31:0] local_bb2_xor_i1640;

assign local_bb2_xor_i1640_inputs_ready = (rnode_169to170_bb2_xor_i1827_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__29_i1856_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_or581_i1885_0_valid_out_1_NO_SHIFT_REG & rnode_169to170_bb2_or581_i1885_0_valid_out_0_NO_SHIFT_REG & rnode_169to170_bb2_reduction_0_i1886_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp68_i1888_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp71_not_i1905_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp77_i1894_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__39_i1897_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and75_i1889_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and74_i1891_0_valid_out_NO_SHIFT_REG);
assign local_bb2_xor_i1640 = (rnode_169to170_bb2__29_i1856_0_NO_SHIFT_REG ? 32'hFFC00000 : local_bb2_or112_i1914_op);
assign local_bb2_xor_i1640_valid_out = 1'b1;
assign rnode_169to170_bb2_xor_i1827_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1856_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i1885_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i1885_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1886_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp68_i1888_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i1905_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i1894_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i1897_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i1889_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and74_i1891_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i1365_stall_local;
wire [31:0] local_bb2_or112_i1365;

assign local_bb2_or112_i1365 = (local_bb2_and108_i1363 | local_bb2_cond111_i1364);

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i628_valid_out;
wire local_bb2_xor_i628_stall_in;
wire local_bb2_xor_i628_inputs_ready;
wire local_bb2_xor_i628_stall_local;
wire [31:0] local_bb2_xor_i628;

assign local_bb2_xor_i628_inputs_ready = (rnode_169to170_bb2_xor_i730_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__29_i759_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_or581_i788_0_valid_out_1_NO_SHIFT_REG & rnode_169to170_bb2_or581_i788_0_valid_out_0_NO_SHIFT_REG & rnode_169to170_bb2_reduction_0_i789_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp68_i791_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp71_not_i808_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_cmp77_i797_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__39_i800_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and75_i792_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and74_i794_0_valid_out_NO_SHIFT_REG);
assign local_bb2_xor_i628 = (rnode_169to170_bb2__29_i759_0_NO_SHIFT_REG ? 32'hFFC00000 : local_bb2_or112_i817_op);
assign local_bb2_xor_i628_valid_out = 1'b1;
assign rnode_169to170_bb2_xor_i730_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i759_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i788_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_or581_i788_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i789_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp68_i791_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp71_not_i808_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i797_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i800_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i792_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and74_i794_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_or112_i353_stall_local;
wire [31:0] local_bb2_or112_i353;

assign local_bb2_or112_i353 = (local_bb2_and108_i351 | local_bb2_cond111_i352);

// This section implements an unregistered operation.
// 
wire local_bb2_and2_i1643_stall_local;
wire [31:0] local_bb2_and2_i1643;

assign local_bb2_and2_i1643 = (rnode_170to171_bb2_var__u94_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and12_i1648_stall_local;
wire [31:0] local_bb2_and12_i1648;

assign local_bb2_and12_i1648 = (rnode_170to171_bb2_var__u94_1_NO_SHIFT_REG & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u95_valid_out;
wire local_bb2_var__u95_stall_in;
wire local_bb2_var__u95_inputs_ready;
wire local_bb2_var__u95_stall_local;
wire [31:0] local_bb2_var__u95;

assign local_bb2_var__u95_inputs_ready = (rnode_169to170_bb2_xor_i1370_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__29_i1399_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_reduction_0_i1429_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_var__u48_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__37_i1426_0_valid_out_0_NO_SHIFT_REG & rnode_169to170_bb2__37_i1426_0_valid_out_1_NO_SHIFT_REG & rnode_169to170_bb2__37_i1426_0_valid_out_3_NO_SHIFT_REG & rnode_169to170_bb2__37_i1426_0_valid_out_2_NO_SHIFT_REG & rnode_169to170_bb2_cmp77_i1437_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__39_i1440_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and75_i1432_0_valid_out_NO_SHIFT_REG);
assign local_bb2_var__u95 = (rnode_169to170_bb2__29_i1399_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb2_or112_i1457);
assign local_bb2_var__u95_valid_out = 1'b1;
assign rnode_169to170_bb2_xor_i1370_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1399_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1429_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u48_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1426_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1426_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1426_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1426_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i1437_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i1440_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i1432_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u96_valid_out;
wire local_bb2_var__u96_stall_in;
wire local_bb2_var__u96_inputs_ready;
wire local_bb2_var__u96_stall_local;
wire [31:0] local_bb2_var__u96;

assign local_bb2_var__u96_inputs_ready = (rnode_169to170_bb2_xor_i822_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__29_i851_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_reduction_0_i881_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_var__u50_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__37_i878_0_valid_out_0_NO_SHIFT_REG & rnode_169to170_bb2__37_i878_0_valid_out_1_NO_SHIFT_REG & rnode_169to170_bb2__37_i878_0_valid_out_3_NO_SHIFT_REG & rnode_169to170_bb2__37_i878_0_valid_out_2_NO_SHIFT_REG & rnode_169to170_bb2_cmp77_i889_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__39_i892_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and75_i884_0_valid_out_NO_SHIFT_REG);
assign local_bb2_var__u96 = (rnode_169to170_bb2__29_i851_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb2_or112_i909);
assign local_bb2_var__u96_valid_out = 1'b1;
assign rnode_169to170_bb2_xor_i822_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i851_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i881_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u50_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i878_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i878_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i878_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i878_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i889_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i892_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i884_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u97_valid_out;
wire local_bb2_var__u97_stall_in;
wire local_bb2_var__u97_inputs_ready;
wire local_bb2_var__u97_stall_local;
wire [31:0] local_bb2_var__u97;

assign local_bb2_var__u97_inputs_ready = (rnode_169to170_bb2_xor_i358_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__29_i387_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_reduction_0_i417_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_var__u52_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__37_i414_0_valid_out_0_NO_SHIFT_REG & rnode_169to170_bb2__37_i414_0_valid_out_1_NO_SHIFT_REG & rnode_169to170_bb2__37_i414_0_valid_out_3_NO_SHIFT_REG & rnode_169to170_bb2__37_i414_0_valid_out_2_NO_SHIFT_REG & rnode_169to170_bb2_cmp77_i425_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__39_i428_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and75_i420_0_valid_out_NO_SHIFT_REG);
assign local_bb2_var__u97 = (rnode_169to170_bb2__29_i387_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb2_or112_i445);
assign local_bb2_var__u97_valid_out = 1'b1;
assign rnode_169to170_bb2_xor_i358_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i387_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i417_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u52_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i414_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i414_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i414_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i414_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i425_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i428_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i420_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb2_xor_i1640_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i1640_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i1640_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i1640_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i1640_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i1640_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i1640_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb2_xor_i1640_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb2_xor_i1640_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb2_xor_i1640_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb2_xor_i1640_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb2_xor_i1640_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i1640),
	.data_out(rnode_170to171_bb2_xor_i1640_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb2_xor_i1640_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_bb2_xor_i1640_0_reg_171_fifo.DATA_WIDTH = 32;
defparam rnode_170to171_bb2_xor_i1640_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_bb2_xor_i1640_0_reg_171_fifo.IMPL = "shift_reg";

assign rnode_170to171_bb2_xor_i1640_0_reg_171_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i1640_stall_in = 1'b0;
assign rnode_170to171_bb2_xor_i1640_0_stall_in_0_reg_171_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i1640_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_xor_i1640_0_NO_SHIFT_REG = rnode_170to171_bb2_xor_i1640_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_xor_i1640_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_xor_i1640_1_NO_SHIFT_REG = rnode_170to171_bb2_xor_i1640_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_xor_i1640_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_xor_i1640_2_NO_SHIFT_REG = rnode_170to171_bb2_xor_i1640_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_xor_i1640_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_xor_i1640_3_NO_SHIFT_REG = rnode_170to171_bb2_xor_i1640_0_reg_171_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u98_valid_out;
wire local_bb2_var__u98_stall_in;
wire local_bb2_var__u98_inputs_ready;
wire local_bb2_var__u98_stall_local;
wire [31:0] local_bb2_var__u98;

assign local_bb2_var__u98_inputs_ready = (rnode_169to170_bb2_xor_i1278_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__29_i1307_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_reduction_0_i1337_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_var__u56_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__37_i1334_0_valid_out_0_NO_SHIFT_REG & rnode_169to170_bb2__37_i1334_0_valid_out_1_NO_SHIFT_REG & rnode_169to170_bb2__37_i1334_0_valid_out_3_NO_SHIFT_REG & rnode_169to170_bb2__37_i1334_0_valid_out_2_NO_SHIFT_REG & rnode_169to170_bb2_cmp77_i1345_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__39_i1348_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and75_i1340_0_valid_out_NO_SHIFT_REG);
assign local_bb2_var__u98 = (rnode_169to170_bb2__29_i1307_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb2_or112_i1365);
assign local_bb2_var__u98_valid_out = 1'b1;
assign rnode_169to170_bb2_xor_i1278_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i1307_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i1337_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u56_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1334_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1334_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1334_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i1334_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i1345_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i1348_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i1340_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb2_xor_i628_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i628_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i628_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i628_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i628_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_xor_i628_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_xor_i628_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb2_xor_i628_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb2_xor_i628_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb2_xor_i628_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb2_xor_i628_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb2_xor_i628_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb2_xor_i628),
	.data_out(rnode_170to171_bb2_xor_i628_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb2_xor_i628_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_bb2_xor_i628_0_reg_171_fifo.DATA_WIDTH = 32;
defparam rnode_170to171_bb2_xor_i628_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_bb2_xor_i628_0_reg_171_fifo.IMPL = "shift_reg";

assign rnode_170to171_bb2_xor_i628_0_reg_171_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_xor_i628_stall_in = 1'b0;
assign rnode_170to171_bb2_xor_i628_0_stall_in_0_reg_171_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i628_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_xor_i628_0_NO_SHIFT_REG = rnode_170to171_bb2_xor_i628_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_xor_i628_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_xor_i628_1_NO_SHIFT_REG = rnode_170to171_bb2_xor_i628_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_xor_i628_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_xor_i628_2_NO_SHIFT_REG = rnode_170to171_bb2_xor_i628_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_xor_i628_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_xor_i628_3_NO_SHIFT_REG = rnode_170to171_bb2_xor_i628_0_reg_171_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u99_valid_out;
wire local_bb2_var__u99_stall_in;
wire local_bb2_var__u99_inputs_ready;
wire local_bb2_var__u99_stall_local;
wire [31:0] local_bb2_var__u99;

assign local_bb2_var__u99_inputs_ready = (rnode_169to170_bb2_xor_i266_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__29_i295_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_reduction_0_i325_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_var__u60_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__37_i322_0_valid_out_0_NO_SHIFT_REG & rnode_169to170_bb2__37_i322_0_valid_out_1_NO_SHIFT_REG & rnode_169to170_bb2__37_i322_0_valid_out_3_NO_SHIFT_REG & rnode_169to170_bb2__37_i322_0_valid_out_2_NO_SHIFT_REG & rnode_169to170_bb2_cmp77_i333_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2__39_i336_0_valid_out_NO_SHIFT_REG & rnode_169to170_bb2_and75_i328_0_valid_out_NO_SHIFT_REG);
assign local_bb2_var__u99 = (rnode_169to170_bb2__29_i295_0_NO_SHIFT_REG ? 32'h7FC00000 : local_bb2_or112_i353);
assign local_bb2_var__u99_valid_out = 1'b1;
assign rnode_169to170_bb2_xor_i266_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__29_i295_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_reduction_0_i325_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_var__u60_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i322_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i322_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i322_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__37_i322_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_cmp77_i333_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2__39_i336_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_169to170_bb2_and75_i328_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i1644_stall_local;
wire [31:0] local_bb2_shr3_i1644;

assign local_bb2_shr3_i1644 = (local_bb2_and2_i1643 & 32'h7FFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb2_var__u95_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u95_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u95_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u95_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u95_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u95_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u95_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb2_var__u95_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb2_var__u95_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb2_var__u95_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb2_var__u95_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb2_var__u95_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb2_var__u95),
	.data_out(rnode_170to171_bb2_var__u95_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb2_var__u95_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_bb2_var__u95_0_reg_171_fifo.DATA_WIDTH = 32;
defparam rnode_170to171_bb2_var__u95_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_bb2_var__u95_0_reg_171_fifo.IMPL = "shift_reg";

assign rnode_170to171_bb2_var__u95_0_reg_171_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u95_stall_in = 1'b0;
assign rnode_170to171_bb2_var__u95_0_stall_in_0_reg_171_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u95_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u95_0_NO_SHIFT_REG = rnode_170to171_bb2_var__u95_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u95_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u95_1_NO_SHIFT_REG = rnode_170to171_bb2_var__u95_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u95_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u95_2_NO_SHIFT_REG = rnode_170to171_bb2_var__u95_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u95_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u95_3_NO_SHIFT_REG = rnode_170to171_bb2_var__u95_0_reg_171_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb2_var__u96_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u96_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u96_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u96_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u96_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u96_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u96_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb2_var__u96_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb2_var__u96_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb2_var__u96_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb2_var__u96_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb2_var__u96_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb2_var__u96),
	.data_out(rnode_170to171_bb2_var__u96_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb2_var__u96_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_bb2_var__u96_0_reg_171_fifo.DATA_WIDTH = 32;
defparam rnode_170to171_bb2_var__u96_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_bb2_var__u96_0_reg_171_fifo.IMPL = "shift_reg";

assign rnode_170to171_bb2_var__u96_0_reg_171_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u96_stall_in = 1'b0;
assign rnode_170to171_bb2_var__u96_0_stall_in_0_reg_171_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u96_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u96_0_NO_SHIFT_REG = rnode_170to171_bb2_var__u96_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u96_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u96_1_NO_SHIFT_REG = rnode_170to171_bb2_var__u96_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u96_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u96_2_NO_SHIFT_REG = rnode_170to171_bb2_var__u96_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u96_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u96_3_NO_SHIFT_REG = rnode_170to171_bb2_var__u96_0_reg_171_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb2_var__u97_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u97_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u97_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u97_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u97_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u97_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u97_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb2_var__u97_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb2_var__u97_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb2_var__u97_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb2_var__u97_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb2_var__u97_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb2_var__u97),
	.data_out(rnode_170to171_bb2_var__u97_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb2_var__u97_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_bb2_var__u97_0_reg_171_fifo.DATA_WIDTH = 32;
defparam rnode_170to171_bb2_var__u97_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_bb2_var__u97_0_reg_171_fifo.IMPL = "shift_reg";

assign rnode_170to171_bb2_var__u97_0_reg_171_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u97_stall_in = 1'b0;
assign rnode_170to171_bb2_var__u97_0_stall_in_0_reg_171_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u97_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u97_0_NO_SHIFT_REG = rnode_170to171_bb2_var__u97_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u97_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u97_1_NO_SHIFT_REG = rnode_170to171_bb2_var__u97_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u97_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u97_2_NO_SHIFT_REG = rnode_170to171_bb2_var__u97_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u97_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u97_3_NO_SHIFT_REG = rnode_170to171_bb2_var__u97_0_reg_171_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and_i1641_stall_local;
wire [31:0] local_bb2_and_i1641;

assign local_bb2_and_i1641 = (rnode_170to171_bb2_xor_i1640_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and10_i1647_stall_local;
wire [31:0] local_bb2_and10_i1647;

assign local_bb2_and10_i1647 = (rnode_170to171_bb2_xor_i1640_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb2_var__u98_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u98_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u98_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u98_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u98_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u98_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u98_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb2_var__u98_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb2_var__u98_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb2_var__u98_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb2_var__u98_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb2_var__u98_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb2_var__u98),
	.data_out(rnode_170to171_bb2_var__u98_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb2_var__u98_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_bb2_var__u98_0_reg_171_fifo.DATA_WIDTH = 32;
defparam rnode_170to171_bb2_var__u98_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_bb2_var__u98_0_reg_171_fifo.IMPL = "shift_reg";

assign rnode_170to171_bb2_var__u98_0_reg_171_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u98_stall_in = 1'b0;
assign rnode_170to171_bb2_var__u98_0_stall_in_0_reg_171_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u98_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u98_0_NO_SHIFT_REG = rnode_170to171_bb2_var__u98_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u98_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u98_1_NO_SHIFT_REG = rnode_170to171_bb2_var__u98_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u98_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u98_2_NO_SHIFT_REG = rnode_170to171_bb2_var__u98_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u98_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u98_3_NO_SHIFT_REG = rnode_170to171_bb2_var__u98_0_reg_171_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and_i629_stall_local;
wire [31:0] local_bb2_and_i629;

assign local_bb2_and_i629 = (rnode_170to171_bb2_xor_i628_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and10_i635_stall_local;
wire [31:0] local_bb2_and10_i635;

assign local_bb2_and10_i635 = (rnode_170to171_bb2_xor_i628_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_170to171_bb2_var__u99_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u99_0_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u99_1_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u99_2_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u99_3_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_reg_171_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_170to171_bb2_var__u99_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_valid_out_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_stall_in_0_reg_171_NO_SHIFT_REG;
 logic rnode_170to171_bb2_var__u99_0_stall_out_reg_171_NO_SHIFT_REG;

acl_data_fifo rnode_170to171_bb2_var__u99_0_reg_171_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_170to171_bb2_var__u99_0_reg_171_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_170to171_bb2_var__u99_0_stall_in_0_reg_171_NO_SHIFT_REG),
	.valid_out(rnode_170to171_bb2_var__u99_0_valid_out_0_reg_171_NO_SHIFT_REG),
	.stall_out(rnode_170to171_bb2_var__u99_0_stall_out_reg_171_NO_SHIFT_REG),
	.data_in(local_bb2_var__u99),
	.data_out(rnode_170to171_bb2_var__u99_0_reg_171_NO_SHIFT_REG)
);

defparam rnode_170to171_bb2_var__u99_0_reg_171_fifo.DEPTH = 1;
defparam rnode_170to171_bb2_var__u99_0_reg_171_fifo.DATA_WIDTH = 32;
defparam rnode_170to171_bb2_var__u99_0_reg_171_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_170to171_bb2_var__u99_0_reg_171_fifo.IMPL = "shift_reg";

assign rnode_170to171_bb2_var__u99_0_reg_171_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u99_stall_in = 1'b0;
assign rnode_170to171_bb2_var__u99_0_stall_in_0_reg_171_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u99_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u99_0_NO_SHIFT_REG = rnode_170to171_bb2_var__u99_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u99_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u99_1_NO_SHIFT_REG = rnode_170to171_bb2_var__u99_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u99_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u99_2_NO_SHIFT_REG = rnode_170to171_bb2_var__u99_0_reg_171_NO_SHIFT_REG;
assign rnode_170to171_bb2_var__u99_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_170to171_bb2_var__u99_3_NO_SHIFT_REG = rnode_170to171_bb2_var__u99_0_reg_171_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and2_i1094_stall_local;
wire [31:0] local_bb2_and2_i1094;

assign local_bb2_and2_i1094 = (rnode_170to171_bb2_var__u95_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and12_i1099_stall_local;
wire [31:0] local_bb2_and12_i1099;

assign local_bb2_and12_i1099 = (rnode_170to171_bb2_var__u95_1_NO_SHIFT_REG & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and2_i631_stall_local;
wire [31:0] local_bb2_and2_i631;

assign local_bb2_and2_i631 = (rnode_170to171_bb2_var__u96_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and12_i636_stall_local;
wire [31:0] local_bb2_and12_i636;

assign local_bb2_and12_i636 = (rnode_170to171_bb2_var__u96_1_NO_SHIFT_REG & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and2_i82_stall_local;
wire [31:0] local_bb2_and2_i82;

assign local_bb2_and2_i82 = (rnode_170to171_bb2_var__u97_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and12_i87_stall_local;
wire [31:0] local_bb2_and12_i87;

assign local_bb2_and12_i87 = (rnode_170to171_bb2_var__u97_1_NO_SHIFT_REG & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i1642_stall_local;
wire [31:0] local_bb2_shr_i1642;

assign local_bb2_shr_i1642 = (local_bb2_and_i1641 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp13_i1649_stall_local;
wire local_bb2_cmp13_i1649;

assign local_bb2_cmp13_i1649 = (local_bb2_and10_i1647 > local_bb2_and12_i1648);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i1092_stall_local;
wire [31:0] local_bb2_and_i1092;

assign local_bb2_and_i1092 = (rnode_170to171_bb2_var__u98_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and10_i1098_stall_local;
wire [31:0] local_bb2_and10_i1098;

assign local_bb2_and10_i1098 = (rnode_170to171_bb2_var__u98_1_NO_SHIFT_REG & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i630_stall_local;
wire [31:0] local_bb2_shr_i630;

assign local_bb2_shr_i630 = (local_bb2_and_i629 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i80_stall_local;
wire [31:0] local_bb2_and_i80;

assign local_bb2_and_i80 = (rnode_170to171_bb2_var__u99_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and10_i86_stall_local;
wire [31:0] local_bb2_and10_i86;

assign local_bb2_and10_i86 = (rnode_170to171_bb2_var__u99_1_NO_SHIFT_REG & 32'hFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i1095_stall_local;
wire [31:0] local_bb2_shr3_i1095;

assign local_bb2_shr3_i1095 = (local_bb2_and2_i1094 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i632_stall_local;
wire [31:0] local_bb2_shr3_i632;

assign local_bb2_shr3_i632 = (local_bb2_and2_i631 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp13_i637_stall_local;
wire local_bb2_cmp13_i637;

assign local_bb2_cmp13_i637 = (local_bb2_and10_i635 > local_bb2_and12_i636);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i83_stall_local;
wire [31:0] local_bb2_shr3_i83;

assign local_bb2_shr3_i83 = (local_bb2_and2_i82 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i1645_stall_local;
wire local_bb2_cmp_i1645;

assign local_bb2_cmp_i1645 = (local_bb2_shr_i1642 > local_bb2_shr3_i1644);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp8_i1646_stall_local;
wire local_bb2_cmp8_i1646;

assign local_bb2_cmp8_i1646 = (local_bb2_shr_i1642 == local_bb2_shr3_i1644);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i1093_stall_local;
wire [31:0] local_bb2_shr_i1093;

assign local_bb2_shr_i1093 = (local_bb2_and_i1092 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp13_i1100_stall_local;
wire local_bb2_cmp13_i1100;

assign local_bb2_cmp13_i1100 = (local_bb2_and10_i1098 > local_bb2_and12_i1099);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i81_stall_local;
wire [31:0] local_bb2_shr_i81;

assign local_bb2_shr_i81 = (local_bb2_and_i80 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp13_i88_stall_local;
wire local_bb2_cmp13_i88;

assign local_bb2_cmp13_i88 = (local_bb2_and10_i86 > local_bb2_and12_i87);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i633_stall_local;
wire local_bb2_cmp_i633;

assign local_bb2_cmp_i633 = (local_bb2_shr_i630 > local_bb2_shr3_i632);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp8_i634_stall_local;
wire local_bb2_cmp8_i634;

assign local_bb2_cmp8_i634 = (local_bb2_shr_i630 == local_bb2_shr3_i632);

// This section implements an unregistered operation.
// 
wire local_bb2___i1650_stall_local;
wire local_bb2___i1650;

assign local_bb2___i1650 = (local_bb2_cmp8_i1646 & local_bb2_cmp13_i1649);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i1096_stall_local;
wire local_bb2_cmp_i1096;

assign local_bb2_cmp_i1096 = (local_bb2_shr_i1093 > local_bb2_shr3_i1095);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp8_i1097_stall_local;
wire local_bb2_cmp8_i1097;

assign local_bb2_cmp8_i1097 = (local_bb2_shr_i1093 == local_bb2_shr3_i1095);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i84_stall_local;
wire local_bb2_cmp_i84;

assign local_bb2_cmp_i84 = (local_bb2_shr_i81 > local_bb2_shr3_i83);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp8_i85_stall_local;
wire local_bb2_cmp8_i85;

assign local_bb2_cmp8_i85 = (local_bb2_shr_i81 == local_bb2_shr3_i83);

// This section implements an unregistered operation.
// 
wire local_bb2___i638_stall_local;
wire local_bb2___i638;

assign local_bb2___i638 = (local_bb2_cmp8_i634 & local_bb2_cmp13_i637);

// This section implements an unregistered operation.
// 
wire local_bb2__21_i1651_stall_local;
wire local_bb2__21_i1651;

assign local_bb2__21_i1651 = (local_bb2_cmp_i1645 | local_bb2___i1650);

// This section implements an unregistered operation.
// 
wire local_bb2___i1101_stall_local;
wire local_bb2___i1101;

assign local_bb2___i1101 = (local_bb2_cmp8_i1097 & local_bb2_cmp13_i1100);

// This section implements an unregistered operation.
// 
wire local_bb2___i89_stall_local;
wire local_bb2___i89;

assign local_bb2___i89 = (local_bb2_cmp8_i85 & local_bb2_cmp13_i88);

// This section implements an unregistered operation.
// 
wire local_bb2__21_i639_stall_local;
wire local_bb2__21_i639;

assign local_bb2__21_i639 = (local_bb2_cmp_i633 | local_bb2___i638);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i1652_stall_local;
wire [31:0] local_bb2__22_i1652;

assign local_bb2__22_i1652 = (local_bb2__21_i1651 ? rnode_170to171_bb2_var__u94_2_NO_SHIFT_REG : rnode_170to171_bb2_xor_i1640_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i1652_valid_out;
wire local_bb2__22_i1652_stall_in;
 reg local_bb2__22_i1652_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i1653_valid_out;
wire local_bb2__23_i1653_stall_in;
 reg local_bb2__23_i1653_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i1653_inputs_ready;
wire local_bb2__23_i1653_stall_local;
wire [31:0] local_bb2__23_i1653;

assign local_bb2__23_i1653_inputs_ready = (rnode_170to171_bb2_var__u94_0_valid_out_0_NO_SHIFT_REG & rnode_170to171_bb2_var__u94_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_bb2_xor_i1640_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_bb2_xor_i1640_0_valid_out_0_NO_SHIFT_REG & rnode_170to171_bb2_var__u94_0_valid_out_2_NO_SHIFT_REG & rnode_170to171_bb2_xor_i1640_0_valid_out_2_NO_SHIFT_REG & rnode_170to171_bb2_xor_i1640_0_valid_out_3_NO_SHIFT_REG & rnode_170to171_bb2_var__u94_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2__23_i1653 = (local_bb2__21_i1651 ? rnode_170to171_bb2_xor_i1640_3_NO_SHIFT_REG : rnode_170to171_bb2_var__u94_3_NO_SHIFT_REG);
assign local_bb2__22_i1652_valid_out = 1'b1;
assign local_bb2__23_i1653_valid_out = 1'b1;
assign rnode_170to171_bb2_var__u94_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u94_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i1640_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i1640_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u94_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i1640_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i1640_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u94_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__22_i1652_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__23_i1653_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__22_i1652_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i1653_inputs_ready & (local_bb2__22_i1652_consumed_0_NO_SHIFT_REG | ~(local_bb2__22_i1652_stall_in)) & local_bb2__23_i1653_stall_local);
		local_bb2__23_i1653_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i1653_inputs_ready & (local_bb2__23_i1653_consumed_0_NO_SHIFT_REG | ~(local_bb2__23_i1653_stall_in)) & local_bb2__23_i1653_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2__21_i1102_stall_local;
wire local_bb2__21_i1102;

assign local_bb2__21_i1102 = (local_bb2_cmp_i1096 | local_bb2___i1101);

// This section implements an unregistered operation.
// 
wire local_bb2__21_i90_stall_local;
wire local_bb2__21_i90;

assign local_bb2__21_i90 = (local_bb2_cmp_i84 | local_bb2___i89);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i640_stall_local;
wire [31:0] local_bb2__22_i640;

assign local_bb2__22_i640 = (local_bb2__21_i639 ? rnode_170to171_bb2_var__u96_2_NO_SHIFT_REG : rnode_170to171_bb2_xor_i628_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i640_valid_out;
wire local_bb2__22_i640_stall_in;
 reg local_bb2__22_i640_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i641_valid_out;
wire local_bb2__23_i641_stall_in;
 reg local_bb2__23_i641_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i641_inputs_ready;
wire local_bb2__23_i641_stall_local;
wire [31:0] local_bb2__23_i641;

assign local_bb2__23_i641_inputs_ready = (rnode_170to171_bb2_var__u96_0_valid_out_0_NO_SHIFT_REG & rnode_170to171_bb2_xor_i628_0_valid_out_0_NO_SHIFT_REG & rnode_170to171_bb2_var__u96_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_bb2_xor_i628_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_bb2_var__u96_0_valid_out_2_NO_SHIFT_REG & rnode_170to171_bb2_xor_i628_0_valid_out_2_NO_SHIFT_REG & rnode_170to171_bb2_xor_i628_0_valid_out_3_NO_SHIFT_REG & rnode_170to171_bb2_var__u96_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2__23_i641 = (local_bb2__21_i639 ? rnode_170to171_bb2_xor_i628_3_NO_SHIFT_REG : rnode_170to171_bb2_var__u96_3_NO_SHIFT_REG);
assign local_bb2__22_i640_valid_out = 1'b1;
assign local_bb2__23_i641_valid_out = 1'b1;
assign rnode_170to171_bb2_var__u96_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i628_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u96_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i628_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u96_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i628_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_xor_i628_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u96_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__22_i640_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__23_i641_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__22_i640_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i641_inputs_ready & (local_bb2__22_i640_consumed_0_NO_SHIFT_REG | ~(local_bb2__22_i640_stall_in)) & local_bb2__23_i641_stall_local);
		local_bb2__23_i641_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i641_inputs_ready & (local_bb2__23_i641_consumed_0_NO_SHIFT_REG | ~(local_bb2__23_i641_stall_in)) & local_bb2__23_i641_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_171to172_bb2__22_i1652_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1652_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i1652_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1652_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1652_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i1652_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1652_0_reg_172_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i1652_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1652_0_valid_out_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1652_0_stall_in_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1652_0_stall_out_reg_172_NO_SHIFT_REG;

acl_data_fifo rnode_171to172_bb2__22_i1652_0_reg_172_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to172_bb2__22_i1652_0_reg_172_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to172_bb2__22_i1652_0_stall_in_0_reg_172_NO_SHIFT_REG),
	.valid_out(rnode_171to172_bb2__22_i1652_0_valid_out_0_reg_172_NO_SHIFT_REG),
	.stall_out(rnode_171to172_bb2__22_i1652_0_stall_out_reg_172_NO_SHIFT_REG),
	.data_in(local_bb2__22_i1652),
	.data_out(rnode_171to172_bb2__22_i1652_0_reg_172_NO_SHIFT_REG)
);

defparam rnode_171to172_bb2__22_i1652_0_reg_172_fifo.DEPTH = 1;
defparam rnode_171to172_bb2__22_i1652_0_reg_172_fifo.DATA_WIDTH = 32;
defparam rnode_171to172_bb2__22_i1652_0_reg_172_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_171to172_bb2__22_i1652_0_reg_172_fifo.IMPL = "shift_reg";

assign rnode_171to172_bb2__22_i1652_0_reg_172_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__22_i1652_stall_in = 1'b0;
assign rnode_171to172_bb2__22_i1652_0_stall_in_0_reg_172_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__22_i1652_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i1652_0_NO_SHIFT_REG = rnode_171to172_bb2__22_i1652_0_reg_172_NO_SHIFT_REG;
assign rnode_171to172_bb2__22_i1652_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i1652_1_NO_SHIFT_REG = rnode_171to172_bb2__22_i1652_0_reg_172_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_171to172_bb2__23_i1653_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1653_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i1653_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1653_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1653_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i1653_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1653_0_reg_172_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i1653_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1653_0_valid_out_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1653_0_stall_in_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1653_0_stall_out_reg_172_NO_SHIFT_REG;

acl_data_fifo rnode_171to172_bb2__23_i1653_0_reg_172_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to172_bb2__23_i1653_0_reg_172_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to172_bb2__23_i1653_0_stall_in_0_reg_172_NO_SHIFT_REG),
	.valid_out(rnode_171to172_bb2__23_i1653_0_valid_out_0_reg_172_NO_SHIFT_REG),
	.stall_out(rnode_171to172_bb2__23_i1653_0_stall_out_reg_172_NO_SHIFT_REG),
	.data_in(local_bb2__23_i1653),
	.data_out(rnode_171to172_bb2__23_i1653_0_reg_172_NO_SHIFT_REG)
);

defparam rnode_171to172_bb2__23_i1653_0_reg_172_fifo.DEPTH = 1;
defparam rnode_171to172_bb2__23_i1653_0_reg_172_fifo.DATA_WIDTH = 32;
defparam rnode_171to172_bb2__23_i1653_0_reg_172_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_171to172_bb2__23_i1653_0_reg_172_fifo.IMPL = "shift_reg";

assign rnode_171to172_bb2__23_i1653_0_reg_172_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__23_i1653_stall_in = 1'b0;
assign rnode_171to172_bb2__23_i1653_0_stall_in_0_reg_172_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__23_i1653_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i1653_0_NO_SHIFT_REG = rnode_171to172_bb2__23_i1653_0_reg_172_NO_SHIFT_REG;
assign rnode_171to172_bb2__23_i1653_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i1653_1_NO_SHIFT_REG = rnode_171to172_bb2__23_i1653_0_reg_172_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__22_i1103_stall_local;
wire [31:0] local_bb2__22_i1103;

assign local_bb2__22_i1103 = (local_bb2__21_i1102 ? rnode_170to171_bb2_var__u95_2_NO_SHIFT_REG : rnode_170to171_bb2_var__u98_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i1103_valid_out;
wire local_bb2__22_i1103_stall_in;
 reg local_bb2__22_i1103_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i1104_valid_out;
wire local_bb2__23_i1104_stall_in;
 reg local_bb2__23_i1104_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i1104_inputs_ready;
wire local_bb2__23_i1104_stall_local;
wire [31:0] local_bb2__23_i1104;

assign local_bb2__23_i1104_inputs_ready = (rnode_170to171_bb2_var__u98_0_valid_out_0_NO_SHIFT_REG & rnode_170to171_bb2_var__u95_0_valid_out_0_NO_SHIFT_REG & rnode_170to171_bb2_var__u98_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_bb2_var__u95_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_bb2_var__u95_0_valid_out_2_NO_SHIFT_REG & rnode_170to171_bb2_var__u98_0_valid_out_2_NO_SHIFT_REG & rnode_170to171_bb2_var__u98_0_valid_out_3_NO_SHIFT_REG & rnode_170to171_bb2_var__u95_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2__23_i1104 = (local_bb2__21_i1102 ? rnode_170to171_bb2_var__u98_3_NO_SHIFT_REG : rnode_170to171_bb2_var__u95_3_NO_SHIFT_REG);
assign local_bb2__22_i1103_valid_out = 1'b1;
assign local_bb2__23_i1104_valid_out = 1'b1;
assign rnode_170to171_bb2_var__u98_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u95_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u98_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u95_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u95_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u98_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u98_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u95_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__22_i1103_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__23_i1104_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__22_i1103_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i1104_inputs_ready & (local_bb2__22_i1103_consumed_0_NO_SHIFT_REG | ~(local_bb2__22_i1103_stall_in)) & local_bb2__23_i1104_stall_local);
		local_bb2__23_i1104_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i1104_inputs_ready & (local_bb2__23_i1104_consumed_0_NO_SHIFT_REG | ~(local_bb2__23_i1104_stall_in)) & local_bb2__23_i1104_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2__22_i91_stall_local;
wire [31:0] local_bb2__22_i91;

assign local_bb2__22_i91 = (local_bb2__21_i90 ? rnode_170to171_bb2_var__u97_2_NO_SHIFT_REG : rnode_170to171_bb2_var__u99_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i91_valid_out;
wire local_bb2__22_i91_stall_in;
 reg local_bb2__22_i91_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i92_valid_out;
wire local_bb2__23_i92_stall_in;
 reg local_bb2__23_i92_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i92_inputs_ready;
wire local_bb2__23_i92_stall_local;
wire [31:0] local_bb2__23_i92;

assign local_bb2__23_i92_inputs_ready = (rnode_170to171_bb2_var__u99_0_valid_out_0_NO_SHIFT_REG & rnode_170to171_bb2_var__u97_0_valid_out_0_NO_SHIFT_REG & rnode_170to171_bb2_var__u99_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_bb2_var__u97_0_valid_out_1_NO_SHIFT_REG & rnode_170to171_bb2_var__u97_0_valid_out_2_NO_SHIFT_REG & rnode_170to171_bb2_var__u99_0_valid_out_2_NO_SHIFT_REG & rnode_170to171_bb2_var__u99_0_valid_out_3_NO_SHIFT_REG & rnode_170to171_bb2_var__u97_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2__23_i92 = (local_bb2__21_i90 ? rnode_170to171_bb2_var__u99_3_NO_SHIFT_REG : rnode_170to171_bb2_var__u97_3_NO_SHIFT_REG);
assign local_bb2__22_i91_valid_out = 1'b1;
assign local_bb2__23_i92_valid_out = 1'b1;
assign rnode_170to171_bb2_var__u99_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u97_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u99_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u97_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u97_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u99_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u99_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_170to171_bb2_var__u97_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__22_i91_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__23_i92_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__22_i91_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i92_inputs_ready & (local_bb2__22_i91_consumed_0_NO_SHIFT_REG | ~(local_bb2__22_i91_stall_in)) & local_bb2__23_i92_stall_local);
		local_bb2__23_i92_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i92_inputs_ready & (local_bb2__23_i92_consumed_0_NO_SHIFT_REG | ~(local_bb2__23_i92_stall_in)) & local_bb2__23_i92_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_171to172_bb2__22_i640_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i640_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i640_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i640_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i640_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i640_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i640_0_reg_172_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i640_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i640_0_valid_out_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i640_0_stall_in_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i640_0_stall_out_reg_172_NO_SHIFT_REG;

acl_data_fifo rnode_171to172_bb2__22_i640_0_reg_172_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to172_bb2__22_i640_0_reg_172_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to172_bb2__22_i640_0_stall_in_0_reg_172_NO_SHIFT_REG),
	.valid_out(rnode_171to172_bb2__22_i640_0_valid_out_0_reg_172_NO_SHIFT_REG),
	.stall_out(rnode_171to172_bb2__22_i640_0_stall_out_reg_172_NO_SHIFT_REG),
	.data_in(local_bb2__22_i640),
	.data_out(rnode_171to172_bb2__22_i640_0_reg_172_NO_SHIFT_REG)
);

defparam rnode_171to172_bb2__22_i640_0_reg_172_fifo.DEPTH = 1;
defparam rnode_171to172_bb2__22_i640_0_reg_172_fifo.DATA_WIDTH = 32;
defparam rnode_171to172_bb2__22_i640_0_reg_172_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_171to172_bb2__22_i640_0_reg_172_fifo.IMPL = "shift_reg";

assign rnode_171to172_bb2__22_i640_0_reg_172_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__22_i640_stall_in = 1'b0;
assign rnode_171to172_bb2__22_i640_0_stall_in_0_reg_172_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__22_i640_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i640_0_NO_SHIFT_REG = rnode_171to172_bb2__22_i640_0_reg_172_NO_SHIFT_REG;
assign rnode_171to172_bb2__22_i640_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i640_1_NO_SHIFT_REG = rnode_171to172_bb2__22_i640_0_reg_172_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_171to172_bb2__23_i641_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i641_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i641_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i641_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i641_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i641_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i641_0_reg_172_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i641_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i641_0_valid_out_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i641_0_stall_in_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i641_0_stall_out_reg_172_NO_SHIFT_REG;

acl_data_fifo rnode_171to172_bb2__23_i641_0_reg_172_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to172_bb2__23_i641_0_reg_172_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to172_bb2__23_i641_0_stall_in_0_reg_172_NO_SHIFT_REG),
	.valid_out(rnode_171to172_bb2__23_i641_0_valid_out_0_reg_172_NO_SHIFT_REG),
	.stall_out(rnode_171to172_bb2__23_i641_0_stall_out_reg_172_NO_SHIFT_REG),
	.data_in(local_bb2__23_i641),
	.data_out(rnode_171to172_bb2__23_i641_0_reg_172_NO_SHIFT_REG)
);

defparam rnode_171to172_bb2__23_i641_0_reg_172_fifo.DEPTH = 1;
defparam rnode_171to172_bb2__23_i641_0_reg_172_fifo.DATA_WIDTH = 32;
defparam rnode_171to172_bb2__23_i641_0_reg_172_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_171to172_bb2__23_i641_0_reg_172_fifo.IMPL = "shift_reg";

assign rnode_171to172_bb2__23_i641_0_reg_172_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__23_i641_stall_in = 1'b0;
assign rnode_171to172_bb2__23_i641_0_stall_in_0_reg_172_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__23_i641_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i641_0_NO_SHIFT_REG = rnode_171to172_bb2__23_i641_0_reg_172_NO_SHIFT_REG;
assign rnode_171to172_bb2__23_i641_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i641_1_NO_SHIFT_REG = rnode_171to172_bb2__23_i641_0_reg_172_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr18_i1656_stall_local;
wire [31:0] local_bb2_shr18_i1656;

assign local_bb2_shr18_i1656 = (rnode_171to172_bb2__22_i1652_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2__22_i1652_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1652_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i1652_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1652_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1652_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i1652_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1652_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i1652_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1652_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1652_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1652_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2__22_i1652_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2__22_i1652_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2__22_i1652_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2__22_i1652_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2__22_i1652_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(rnode_171to172_bb2__22_i1652_1_NO_SHIFT_REG),
	.data_out(rnode_172to173_bb2__22_i1652_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2__22_i1652_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2__22_i1652_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2__22_i1652_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2__22_i1652_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2__22_i1652_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i1652_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i1652_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i1652_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__22_i1652_0_NO_SHIFT_REG = rnode_172to173_bb2__22_i1652_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__22_i1652_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__22_i1652_1_NO_SHIFT_REG = rnode_172to173_bb2__22_i1652_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i1654_stall_local;
wire [31:0] local_bb2_shr16_i1654;

assign local_bb2_shr16_i1654 = (rnode_171to172_bb2__23_i1653_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2__23_i1653_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i1653_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i1653_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i1653_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i1653_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1653_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2__23_i1653_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2__23_i1653_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2__23_i1653_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2__23_i1653_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2__23_i1653_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(rnode_171to172_bb2__23_i1653_1_NO_SHIFT_REG),
	.data_out(rnode_172to173_bb2__23_i1653_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2__23_i1653_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2__23_i1653_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2__23_i1653_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2__23_i1653_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2__23_i1653_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i1653_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i1653_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i1653_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i1653_0_NO_SHIFT_REG = rnode_172to173_bb2__23_i1653_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__23_i1653_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i1653_1_NO_SHIFT_REG = rnode_172to173_bb2__23_i1653_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__23_i1653_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i1653_2_NO_SHIFT_REG = rnode_172to173_bb2__23_i1653_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_171to172_bb2__22_i1103_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1103_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i1103_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1103_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1103_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i1103_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1103_0_reg_172_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i1103_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1103_0_valid_out_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1103_0_stall_in_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i1103_0_stall_out_reg_172_NO_SHIFT_REG;

acl_data_fifo rnode_171to172_bb2__22_i1103_0_reg_172_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to172_bb2__22_i1103_0_reg_172_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to172_bb2__22_i1103_0_stall_in_0_reg_172_NO_SHIFT_REG),
	.valid_out(rnode_171to172_bb2__22_i1103_0_valid_out_0_reg_172_NO_SHIFT_REG),
	.stall_out(rnode_171to172_bb2__22_i1103_0_stall_out_reg_172_NO_SHIFT_REG),
	.data_in(local_bb2__22_i1103),
	.data_out(rnode_171to172_bb2__22_i1103_0_reg_172_NO_SHIFT_REG)
);

defparam rnode_171to172_bb2__22_i1103_0_reg_172_fifo.DEPTH = 1;
defparam rnode_171to172_bb2__22_i1103_0_reg_172_fifo.DATA_WIDTH = 32;
defparam rnode_171to172_bb2__22_i1103_0_reg_172_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_171to172_bb2__22_i1103_0_reg_172_fifo.IMPL = "shift_reg";

assign rnode_171to172_bb2__22_i1103_0_reg_172_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__22_i1103_stall_in = 1'b0;
assign rnode_171to172_bb2__22_i1103_0_stall_in_0_reg_172_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__22_i1103_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i1103_0_NO_SHIFT_REG = rnode_171to172_bb2__22_i1103_0_reg_172_NO_SHIFT_REG;
assign rnode_171to172_bb2__22_i1103_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i1103_1_NO_SHIFT_REG = rnode_171to172_bb2__22_i1103_0_reg_172_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_171to172_bb2__23_i1104_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1104_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i1104_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1104_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1104_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i1104_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1104_0_reg_172_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i1104_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1104_0_valid_out_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1104_0_stall_in_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i1104_0_stall_out_reg_172_NO_SHIFT_REG;

acl_data_fifo rnode_171to172_bb2__23_i1104_0_reg_172_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to172_bb2__23_i1104_0_reg_172_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to172_bb2__23_i1104_0_stall_in_0_reg_172_NO_SHIFT_REG),
	.valid_out(rnode_171to172_bb2__23_i1104_0_valid_out_0_reg_172_NO_SHIFT_REG),
	.stall_out(rnode_171to172_bb2__23_i1104_0_stall_out_reg_172_NO_SHIFT_REG),
	.data_in(local_bb2__23_i1104),
	.data_out(rnode_171to172_bb2__23_i1104_0_reg_172_NO_SHIFT_REG)
);

defparam rnode_171to172_bb2__23_i1104_0_reg_172_fifo.DEPTH = 1;
defparam rnode_171to172_bb2__23_i1104_0_reg_172_fifo.DATA_WIDTH = 32;
defparam rnode_171to172_bb2__23_i1104_0_reg_172_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_171to172_bb2__23_i1104_0_reg_172_fifo.IMPL = "shift_reg";

assign rnode_171to172_bb2__23_i1104_0_reg_172_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__23_i1104_stall_in = 1'b0;
assign rnode_171to172_bb2__23_i1104_0_stall_in_0_reg_172_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__23_i1104_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i1104_0_NO_SHIFT_REG = rnode_171to172_bb2__23_i1104_0_reg_172_NO_SHIFT_REG;
assign rnode_171to172_bb2__23_i1104_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i1104_1_NO_SHIFT_REG = rnode_171to172_bb2__23_i1104_0_reg_172_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_171to172_bb2__22_i91_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i91_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i91_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i91_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i91_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i91_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i91_0_reg_172_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__22_i91_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i91_0_valid_out_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i91_0_stall_in_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__22_i91_0_stall_out_reg_172_NO_SHIFT_REG;

acl_data_fifo rnode_171to172_bb2__22_i91_0_reg_172_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to172_bb2__22_i91_0_reg_172_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to172_bb2__22_i91_0_stall_in_0_reg_172_NO_SHIFT_REG),
	.valid_out(rnode_171to172_bb2__22_i91_0_valid_out_0_reg_172_NO_SHIFT_REG),
	.stall_out(rnode_171to172_bb2__22_i91_0_stall_out_reg_172_NO_SHIFT_REG),
	.data_in(local_bb2__22_i91),
	.data_out(rnode_171to172_bb2__22_i91_0_reg_172_NO_SHIFT_REG)
);

defparam rnode_171to172_bb2__22_i91_0_reg_172_fifo.DEPTH = 1;
defparam rnode_171to172_bb2__22_i91_0_reg_172_fifo.DATA_WIDTH = 32;
defparam rnode_171to172_bb2__22_i91_0_reg_172_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_171to172_bb2__22_i91_0_reg_172_fifo.IMPL = "shift_reg";

assign rnode_171to172_bb2__22_i91_0_reg_172_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__22_i91_stall_in = 1'b0;
assign rnode_171to172_bb2__22_i91_0_stall_in_0_reg_172_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__22_i91_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i91_0_NO_SHIFT_REG = rnode_171to172_bb2__22_i91_0_reg_172_NO_SHIFT_REG;
assign rnode_171to172_bb2__22_i91_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i91_1_NO_SHIFT_REG = rnode_171to172_bb2__22_i91_0_reg_172_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_171to172_bb2__23_i92_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i92_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i92_0_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i92_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i92_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i92_1_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i92_0_reg_172_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_171to172_bb2__23_i92_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i92_0_valid_out_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i92_0_stall_in_0_reg_172_NO_SHIFT_REG;
 logic rnode_171to172_bb2__23_i92_0_stall_out_reg_172_NO_SHIFT_REG;

acl_data_fifo rnode_171to172_bb2__23_i92_0_reg_172_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_171to172_bb2__23_i92_0_reg_172_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_171to172_bb2__23_i92_0_stall_in_0_reg_172_NO_SHIFT_REG),
	.valid_out(rnode_171to172_bb2__23_i92_0_valid_out_0_reg_172_NO_SHIFT_REG),
	.stall_out(rnode_171to172_bb2__23_i92_0_stall_out_reg_172_NO_SHIFT_REG),
	.data_in(local_bb2__23_i92),
	.data_out(rnode_171to172_bb2__23_i92_0_reg_172_NO_SHIFT_REG)
);

defparam rnode_171to172_bb2__23_i92_0_reg_172_fifo.DEPTH = 1;
defparam rnode_171to172_bb2__23_i92_0_reg_172_fifo.DATA_WIDTH = 32;
defparam rnode_171to172_bb2__23_i92_0_reg_172_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_171to172_bb2__23_i92_0_reg_172_fifo.IMPL = "shift_reg";

assign rnode_171to172_bb2__23_i92_0_reg_172_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__23_i92_stall_in = 1'b0;
assign rnode_171to172_bb2__23_i92_0_stall_in_0_reg_172_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__23_i92_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i92_0_NO_SHIFT_REG = rnode_171to172_bb2__23_i92_0_reg_172_NO_SHIFT_REG;
assign rnode_171to172_bb2__23_i92_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i92_1_NO_SHIFT_REG = rnode_171to172_bb2__23_i92_0_reg_172_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr18_i644_stall_local;
wire [31:0] local_bb2_shr18_i644;

assign local_bb2_shr18_i644 = (rnode_171to172_bb2__22_i640_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2__22_i640_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i640_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i640_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i640_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i640_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i640_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i640_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i640_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i640_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i640_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i640_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2__22_i640_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2__22_i640_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2__22_i640_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2__22_i640_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2__22_i640_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(rnode_171to172_bb2__22_i640_1_NO_SHIFT_REG),
	.data_out(rnode_172to173_bb2__22_i640_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2__22_i640_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2__22_i640_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2__22_i640_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2__22_i640_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2__22_i640_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i640_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i640_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i640_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__22_i640_0_NO_SHIFT_REG = rnode_172to173_bb2__22_i640_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__22_i640_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__22_i640_1_NO_SHIFT_REG = rnode_172to173_bb2__22_i640_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i642_stall_local;
wire [31:0] local_bb2_shr16_i642;

assign local_bb2_shr16_i642 = (rnode_171to172_bb2__23_i641_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2__23_i641_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i641_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i641_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i641_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i641_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i641_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2__23_i641_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2__23_i641_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2__23_i641_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2__23_i641_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2__23_i641_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(rnode_171to172_bb2__23_i641_1_NO_SHIFT_REG),
	.data_out(rnode_172to173_bb2__23_i641_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2__23_i641_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2__23_i641_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2__23_i641_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2__23_i641_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2__23_i641_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i641_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i641_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i641_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i641_0_NO_SHIFT_REG = rnode_172to173_bb2__23_i641_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__23_i641_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i641_1_NO_SHIFT_REG = rnode_172to173_bb2__23_i641_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__23_i641_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i641_2_NO_SHIFT_REG = rnode_172to173_bb2__23_i641_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and19_i1657_stall_local;
wire [31:0] local_bb2_and19_i1657;

assign local_bb2_and19_i1657 = (local_bb2_shr18_i1656 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and21_i1659_stall_local;
wire [31:0] local_bb2_and21_i1659;

assign local_bb2_and21_i1659 = (rnode_172to173_bb2__22_i1652_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i1686_stall_local;
wire [31:0] local_bb2_sub_i1686;

assign local_bb2_sub_i1686 = (local_bb2_shr16_i1654 - local_bb2_shr18_i1656);

// This section implements an unregistered operation.
// 
wire local_bb2_and20_i1658_stall_local;
wire [31:0] local_bb2_and20_i1658;

assign local_bb2_and20_i1658 = (rnode_172to173_bb2__23_i1653_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and35_i1664_valid_out;
wire local_bb2_and35_i1664_stall_in;
wire local_bb2_and35_i1664_inputs_ready;
wire local_bb2_and35_i1664_stall_local;
wire [31:0] local_bb2_and35_i1664;

assign local_bb2_and35_i1664_inputs_ready = rnode_172to173_bb2__23_i1653_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and35_i1664 = (rnode_172to173_bb2__23_i1653_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb2_and35_i1664_valid_out = 1'b1;
assign rnode_172to173_bb2__23_i1653_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_xor36_i1665_stall_local;
wire [31:0] local_bb2_xor36_i1665;

assign local_bb2_xor36_i1665 = (rnode_172to173_bb2__23_i1653_2_NO_SHIFT_REG ^ rnode_172to173_bb2__22_i1652_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shr18_i1107_stall_local;
wire [31:0] local_bb2_shr18_i1107;

assign local_bb2_shr18_i1107 = (rnode_171to172_bb2__22_i1103_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2__22_i1103_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1103_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i1103_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1103_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1103_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i1103_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1103_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i1103_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1103_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1103_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i1103_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2__22_i1103_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2__22_i1103_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2__22_i1103_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2__22_i1103_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2__22_i1103_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(rnode_171to172_bb2__22_i1103_1_NO_SHIFT_REG),
	.data_out(rnode_172to173_bb2__22_i1103_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2__22_i1103_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2__22_i1103_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2__22_i1103_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2__22_i1103_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2__22_i1103_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i1103_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i1103_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i1103_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__22_i1103_0_NO_SHIFT_REG = rnode_172to173_bb2__22_i1103_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__22_i1103_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__22_i1103_1_NO_SHIFT_REG = rnode_172to173_bb2__22_i1103_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i1105_stall_local;
wire [31:0] local_bb2_shr16_i1105;

assign local_bb2_shr16_i1105 = (rnode_171to172_bb2__23_i1104_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2__23_i1104_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i1104_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i1104_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i1104_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i1104_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i1104_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2__23_i1104_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2__23_i1104_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2__23_i1104_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2__23_i1104_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2__23_i1104_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(rnode_171to172_bb2__23_i1104_1_NO_SHIFT_REG),
	.data_out(rnode_172to173_bb2__23_i1104_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2__23_i1104_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2__23_i1104_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2__23_i1104_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2__23_i1104_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2__23_i1104_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i1104_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i1104_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i1104_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i1104_0_NO_SHIFT_REG = rnode_172to173_bb2__23_i1104_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__23_i1104_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i1104_1_NO_SHIFT_REG = rnode_172to173_bb2__23_i1104_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__23_i1104_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i1104_2_NO_SHIFT_REG = rnode_172to173_bb2__23_i1104_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr18_i95_stall_local;
wire [31:0] local_bb2_shr18_i95;

assign local_bb2_shr18_i95 = (rnode_171to172_bb2__22_i91_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2__22_i91_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i91_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i91_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i91_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i91_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i91_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i91_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__22_i91_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i91_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i91_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__22_i91_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2__22_i91_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2__22_i91_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2__22_i91_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2__22_i91_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2__22_i91_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(rnode_171to172_bb2__22_i91_1_NO_SHIFT_REG),
	.data_out(rnode_172to173_bb2__22_i91_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2__22_i91_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2__22_i91_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2__22_i91_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2__22_i91_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2__22_i91_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__22_i91_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i91_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i91_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__22_i91_0_NO_SHIFT_REG = rnode_172to173_bb2__22_i91_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__22_i91_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__22_i91_1_NO_SHIFT_REG = rnode_172to173_bb2__22_i91_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i93_stall_local;
wire [31:0] local_bb2_shr16_i93;

assign local_bb2_shr16_i93 = (rnode_171to172_bb2__23_i92_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2__23_i92_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i92_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i92_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i92_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2__23_i92_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2__23_i92_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2__23_i92_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2__23_i92_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2__23_i92_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2__23_i92_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2__23_i92_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(rnode_171to172_bb2__23_i92_1_NO_SHIFT_REG),
	.data_out(rnode_172to173_bb2__23_i92_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2__23_i92_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2__23_i92_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2__23_i92_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2__23_i92_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2__23_i92_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_171to172_bb2__23_i92_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i92_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i92_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i92_0_NO_SHIFT_REG = rnode_172to173_bb2__23_i92_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__23_i92_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i92_1_NO_SHIFT_REG = rnode_172to173_bb2__23_i92_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2__23_i92_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2__23_i92_2_NO_SHIFT_REG = rnode_172to173_bb2__23_i92_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and19_i645_stall_local;
wire [31:0] local_bb2_and19_i645;

assign local_bb2_and19_i645 = (local_bb2_shr18_i644 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and21_i647_stall_local;
wire [31:0] local_bb2_and21_i647;

assign local_bb2_and21_i647 = (rnode_172to173_bb2__22_i640_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i670_stall_local;
wire [31:0] local_bb2_sub_i670;

assign local_bb2_sub_i670 = (local_bb2_shr16_i642 - local_bb2_shr18_i644);

// This section implements an unregistered operation.
// 
wire local_bb2_and20_i646_stall_local;
wire [31:0] local_bb2_and20_i646;

assign local_bb2_and20_i646 = (rnode_172to173_bb2__23_i641_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and35_i652_valid_out;
wire local_bb2_and35_i652_stall_in;
wire local_bb2_and35_i652_inputs_ready;
wire local_bb2_and35_i652_stall_local;
wire [31:0] local_bb2_and35_i652;

assign local_bb2_and35_i652_inputs_ready = rnode_172to173_bb2__23_i641_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and35_i652 = (rnode_172to173_bb2__23_i641_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb2_and35_i652_valid_out = 1'b1;
assign rnode_172to173_bb2__23_i641_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_xor36_i_stall_local;
wire [31:0] local_bb2_xor36_i;

assign local_bb2_xor36_i = (rnode_172to173_bb2__23_i641_2_NO_SHIFT_REG ^ rnode_172to173_bb2__22_i640_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot23_i1661_stall_local;
wire local_bb2_lnot23_i1661;

assign local_bb2_lnot23_i1661 = (local_bb2_and19_i1657 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp27_i1663_stall_local;
wire local_bb2_cmp27_i1663;

assign local_bb2_cmp27_i1663 = (local_bb2_and19_i1657 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot33_not_i1670_stall_local;
wire local_bb2_lnot33_not_i1670;

assign local_bb2_lnot33_not_i1670 = (local_bb2_and21_i1659 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or65_i1683_stall_local;
wire [31:0] local_bb2_or65_i1683;

assign local_bb2_or65_i1683 = (local_bb2_and21_i1659 << 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and69_i1687_stall_local;
wire [31:0] local_bb2_and69_i1687;

assign local_bb2_and69_i1687 = (local_bb2_sub_i1686 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_i1668_stall_local;
wire local_bb2_lnot30_i1668;

assign local_bb2_lnot30_i1668 = (local_bb2_and20_i1658 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i1680_stall_local;
wire [31:0] local_bb2_or_i1680;

assign local_bb2_or_i1680 = (local_bb2_and20_i1658 << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_and35_i1664_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1664_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_and35_i1664_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1664_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_and35_i1664_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1664_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1664_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1664_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_and35_i1664_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_and35_i1664_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_and35_i1664_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_and35_i1664_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_and35_i1664_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_and35_i1664),
	.data_out(rnode_173to174_bb2_and35_i1664_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_and35_i1664_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_and35_i1664_0_reg_174_fifo.DATA_WIDTH = 32;
defparam rnode_173to174_bb2_and35_i1664_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_and35_i1664_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_and35_i1664_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and35_i1664_stall_in = 1'b0;
assign rnode_173to174_bb2_and35_i1664_0_NO_SHIFT_REG = rnode_173to174_bb2_and35_i1664_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_and35_i1664_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_and35_i1664_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp38_i1666_stall_local;
wire local_bb2_cmp38_i1666;

assign local_bb2_cmp38_i1666 = ($signed(local_bb2_xor36_i1665) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_xor36_lobit_i1739_stall_local;
wire [31:0] local_bb2_xor36_lobit_i1739;

assign local_bb2_xor36_lobit_i1739 = ($signed(local_bb2_xor36_i1665) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and37_lobit_i1741_stall_local;
wire [31:0] local_bb2_and37_lobit_i1741;

assign local_bb2_and37_lobit_i1741 = (local_bb2_xor36_i1665 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and19_i1108_stall_local;
wire [31:0] local_bb2_and19_i1108;

assign local_bb2_and19_i1108 = (local_bb2_shr18_i1107 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and21_i1110_stall_local;
wire [31:0] local_bb2_and21_i1110;

assign local_bb2_and21_i1110 = (rnode_172to173_bb2__22_i1103_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i1137_stall_local;
wire [31:0] local_bb2_sub_i1137;

assign local_bb2_sub_i1137 = (local_bb2_shr16_i1105 - local_bb2_shr18_i1107);

// This section implements an unregistered operation.
// 
wire local_bb2_and20_i1109_stall_local;
wire [31:0] local_bb2_and20_i1109;

assign local_bb2_and20_i1109 = (rnode_172to173_bb2__23_i1104_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and35_i1115_valid_out;
wire local_bb2_and35_i1115_stall_in;
wire local_bb2_and35_i1115_inputs_ready;
wire local_bb2_and35_i1115_stall_local;
wire [31:0] local_bb2_and35_i1115;

assign local_bb2_and35_i1115_inputs_ready = rnode_172to173_bb2__23_i1104_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and35_i1115 = (rnode_172to173_bb2__23_i1104_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb2_and35_i1115_valid_out = 1'b1;
assign rnode_172to173_bb2__23_i1104_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i1116_stall_local;
wire [31:0] local_bb2_xor_i1116;

assign local_bb2_xor_i1116 = (rnode_172to173_bb2__23_i1104_2_NO_SHIFT_REG ^ rnode_172to173_bb2__22_i1103_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and19_i96_stall_local;
wire [31:0] local_bb2_and19_i96;

assign local_bb2_and19_i96 = (local_bb2_shr18_i95 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and21_i98_stall_local;
wire [31:0] local_bb2_and21_i98;

assign local_bb2_and21_i98 = (rnode_172to173_bb2__22_i91_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i125_stall_local;
wire [31:0] local_bb2_sub_i125;

assign local_bb2_sub_i125 = (local_bb2_shr16_i93 - local_bb2_shr18_i95);

// This section implements an unregistered operation.
// 
wire local_bb2_and20_i97_stall_local;
wire [31:0] local_bb2_and20_i97;

assign local_bb2_and20_i97 = (rnode_172to173_bb2__23_i92_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and35_i103_valid_out;
wire local_bb2_and35_i103_stall_in;
wire local_bb2_and35_i103_inputs_ready;
wire local_bb2_and35_i103_stall_local;
wire [31:0] local_bb2_and35_i103;

assign local_bb2_and35_i103_inputs_ready = rnode_172to173_bb2__23_i92_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and35_i103 = (rnode_172to173_bb2__23_i92_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb2_and35_i103_valid_out = 1'b1;
assign rnode_172to173_bb2__23_i92_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i104_stall_local;
wire [31:0] local_bb2_xor_i104;

assign local_bb2_xor_i104 = (rnode_172to173_bb2__23_i92_2_NO_SHIFT_REG ^ rnode_172to173_bb2__22_i91_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot23_i649_stall_local;
wire local_bb2_lnot23_i649;

assign local_bb2_lnot23_i649 = (local_bb2_and19_i645 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp27_i651_stall_local;
wire local_bb2_cmp27_i651;

assign local_bb2_cmp27_i651 = (local_bb2_and19_i645 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot33_not_i656_stall_local;
wire local_bb2_lnot33_not_i656;

assign local_bb2_lnot33_not_i656 = (local_bb2_and21_i647 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or65_i_stall_local;
wire [31:0] local_bb2_or65_i;

assign local_bb2_or65_i = (local_bb2_and21_i647 << 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and69_i_stall_local;
wire [31:0] local_bb2_and69_i;

assign local_bb2_and69_i = (local_bb2_sub_i670 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_i654_stall_local;
wire local_bb2_lnot30_i654;

assign local_bb2_lnot30_i654 = (local_bb2_and20_i646 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i666_stall_local;
wire [31:0] local_bb2_or_i666;

assign local_bb2_or_i666 = (local_bb2_and20_i646 << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_and35_i652_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i652_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_and35_i652_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i652_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_and35_i652_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i652_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i652_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i652_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_and35_i652_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_and35_i652_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_and35_i652_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_and35_i652_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_and35_i652_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_and35_i652),
	.data_out(rnode_173to174_bb2_and35_i652_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_and35_i652_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_and35_i652_0_reg_174_fifo.DATA_WIDTH = 32;
defparam rnode_173to174_bb2_and35_i652_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_and35_i652_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_and35_i652_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and35_i652_stall_in = 1'b0;
assign rnode_173to174_bb2_and35_i652_0_NO_SHIFT_REG = rnode_173to174_bb2_and35_i652_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_and35_i652_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_and35_i652_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp38_i_stall_local;
wire local_bb2_cmp38_i;

assign local_bb2_cmp38_i = ($signed(local_bb2_xor36_i) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_xor36_lobit_i_stall_local;
wire [31:0] local_bb2_xor36_lobit_i;

assign local_bb2_xor36_lobit_i = ($signed(local_bb2_xor36_i) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and37_lobit_i_stall_local;
wire [31:0] local_bb2_and37_lobit_i;

assign local_bb2_and37_lobit_i = (local_bb2_xor36_i >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_shl66_i1684_stall_local;
wire [31:0] local_bb2_shl66_i1684;

assign local_bb2_shl66_i1684 = (local_bb2_or65_i1683 | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp70_i1688_stall_local;
wire local_bb2_cmp70_i1688;

assign local_bb2_cmp70_i1688 = (local_bb2_and69_i1687 > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_not_i1672_stall_local;
wire local_bb2_lnot30_not_i1672;

assign local_bb2_lnot30_not_i1672 = (local_bb2_lnot30_i1668 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i1681_stall_local;
wire [31:0] local_bb2_shl_i1681;

assign local_bb2_shl_i1681 = (local_bb2_or_i1680 | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and35_i1664_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1664_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and35_i1664_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1664_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and35_i1664_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1664_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1664_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1664_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and35_i1664_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and35_i1664_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and35_i1664_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and35_i1664_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and35_i1664_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2_and35_i1664_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2_and35_i1664_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and35_i1664_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and35_i1664_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and35_i1664_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and35_i1664_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and35_i1664_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_and35_i1664_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and35_i1664_0_NO_SHIFT_REG = rnode_174to175_bb2_and35_i1664_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and35_i1664_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and35_i1664_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot23_i1112_stall_local;
wire local_bb2_lnot23_i1112;

assign local_bb2_lnot23_i1112 = (local_bb2_and19_i1108 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp27_i1114_stall_local;
wire local_bb2_cmp27_i1114;

assign local_bb2_cmp27_i1114 = (local_bb2_and19_i1108 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot33_not_i1121_stall_local;
wire local_bb2_lnot33_not_i1121;

assign local_bb2_lnot33_not_i1121 = (local_bb2_and21_i1110 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or64_i1134_stall_local;
wire [31:0] local_bb2_or64_i1134;

assign local_bb2_or64_i1134 = (local_bb2_and21_i1110 << 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and68_i1138_stall_local;
wire [31:0] local_bb2_and68_i1138;

assign local_bb2_and68_i1138 = (local_bb2_sub_i1137 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_i1119_stall_local;
wire local_bb2_lnot30_i1119;

assign local_bb2_lnot30_i1119 = (local_bb2_and20_i1109 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i1131_stall_local;
wire [31:0] local_bb2_or_i1131;

assign local_bb2_or_i1131 = (local_bb2_and20_i1109 << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_and35_i1115_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1115_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_and35_i1115_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1115_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_and35_i1115_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1115_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1115_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i1115_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_and35_i1115_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_and35_i1115_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_and35_i1115_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_and35_i1115_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_and35_i1115_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_and35_i1115),
	.data_out(rnode_173to174_bb2_and35_i1115_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_and35_i1115_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_and35_i1115_0_reg_174_fifo.DATA_WIDTH = 32;
defparam rnode_173to174_bb2_and35_i1115_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_and35_i1115_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_and35_i1115_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and35_i1115_stall_in = 1'b0;
assign rnode_173to174_bb2_and35_i1115_0_NO_SHIFT_REG = rnode_173to174_bb2_and35_i1115_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_and35_i1115_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_and35_i1115_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i1117_stall_local;
wire local_bb2_cmp37_i1117;

assign local_bb2_cmp37_i1117 = ($signed(local_bb2_xor_i1116) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_xor_lobit_i1190_stall_local;
wire [31:0] local_bb2_xor_lobit_i1190;

assign local_bb2_xor_lobit_i1190 = ($signed(local_bb2_xor_i1116) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and36_lobit_i1192_stall_local;
wire [31:0] local_bb2_and36_lobit_i1192;

assign local_bb2_and36_lobit_i1192 = (local_bb2_xor_i1116 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot23_i100_stall_local;
wire local_bb2_lnot23_i100;

assign local_bb2_lnot23_i100 = (local_bb2_and19_i96 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp27_i102_stall_local;
wire local_bb2_cmp27_i102;

assign local_bb2_cmp27_i102 = (local_bb2_and19_i96 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot33_not_i109_stall_local;
wire local_bb2_lnot33_not_i109;

assign local_bb2_lnot33_not_i109 = (local_bb2_and21_i98 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or64_i122_stall_local;
wire [31:0] local_bb2_or64_i122;

assign local_bb2_or64_i122 = (local_bb2_and21_i98 << 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and68_i126_stall_local;
wire [31:0] local_bb2_and68_i126;

assign local_bb2_and68_i126 = (local_bb2_sub_i125 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_i107_stall_local;
wire local_bb2_lnot30_i107;

assign local_bb2_lnot30_i107 = (local_bb2_and20_i97 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i119_stall_local;
wire [31:0] local_bb2_or_i119;

assign local_bb2_or_i119 = (local_bb2_and20_i97 << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_and35_i103_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i103_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_and35_i103_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i103_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_and35_i103_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i103_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i103_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_and35_i103_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_and35_i103_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_and35_i103_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_and35_i103_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_and35_i103_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_and35_i103_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_and35_i103),
	.data_out(rnode_173to174_bb2_and35_i103_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_and35_i103_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_and35_i103_0_reg_174_fifo.DATA_WIDTH = 32;
defparam rnode_173to174_bb2_and35_i103_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_and35_i103_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_and35_i103_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and35_i103_stall_in = 1'b0;
assign rnode_173to174_bb2_and35_i103_0_NO_SHIFT_REG = rnode_173to174_bb2_and35_i103_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_and35_i103_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_and35_i103_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i105_stall_local;
wire local_bb2_cmp37_i105;

assign local_bb2_cmp37_i105 = ($signed(local_bb2_xor_i104) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_xor_lobit_i178_stall_local;
wire [31:0] local_bb2_xor_lobit_i178;

assign local_bb2_xor_lobit_i178 = ($signed(local_bb2_xor_i104) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and36_lobit_i180_stall_local;
wire [31:0] local_bb2_and36_lobit_i180;

assign local_bb2_and36_lobit_i180 = (local_bb2_xor_i104 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_shl66_i_stall_local;
wire [31:0] local_bb2_shl66_i;

assign local_bb2_shl66_i = (local_bb2_or65_i | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp70_i_stall_local;
wire local_bb2_cmp70_i;

assign local_bb2_cmp70_i = (local_bb2_and69_i > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_not_i658_stall_local;
wire local_bb2_lnot30_not_i658;

assign local_bb2_lnot30_not_i658 = (local_bb2_lnot30_i654 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i667_stall_local;
wire [31:0] local_bb2_shl_i667;

assign local_bb2_shl_i667 = (local_bb2_or_i666 | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and35_i652_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i652_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and35_i652_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i652_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and35_i652_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i652_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i652_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i652_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and35_i652_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and35_i652_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and35_i652_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and35_i652_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and35_i652_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2_and35_i652_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2_and35_i652_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and35_i652_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and35_i652_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and35_i652_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and35_i652_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and35_i652_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_and35_i652_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and35_i652_0_NO_SHIFT_REG = rnode_174to175_bb2_and35_i652_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and35_i652_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and35_i652_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i1654_valid_out_1;
wire local_bb2_shr16_i1654_stall_in_1;
 reg local_bb2_shr16_i1654_consumed_1_NO_SHIFT_REG;
wire local_bb2_lnot23_i1661_valid_out;
wire local_bb2_lnot23_i1661_stall_in;
 reg local_bb2_lnot23_i1661_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp27_i1663_valid_out;
wire local_bb2_cmp27_i1663_stall_in;
 reg local_bb2_cmp27_i1663_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i1689_valid_out;
wire local_bb2_align_0_i1689_stall_in;
 reg local_bb2_align_0_i1689_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i1689_inputs_ready;
wire local_bb2_align_0_i1689_stall_local;
wire [31:0] local_bb2_align_0_i1689;

assign local_bb2_align_0_i1689_inputs_ready = (rnode_171to172_bb2__22_i1652_0_valid_out_0_NO_SHIFT_REG & rnode_171to172_bb2__23_i1653_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_align_0_i1689 = (local_bb2_cmp70_i1688 ? 32'h1F : local_bb2_and69_i1687);
assign local_bb2_shr16_i1654_valid_out_1 = 1'b1;
assign local_bb2_lnot23_i1661_valid_out = 1'b1;
assign local_bb2_cmp27_i1663_valid_out = 1'b1;
assign local_bb2_align_0_i1689_valid_out = 1'b1;
assign rnode_171to172_bb2__22_i1652_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__23_i1653_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_shr16_i1654_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lnot23_i1661_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp27_i1663_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_align_0_i1689_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_shr16_i1654_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i1689_inputs_ready & (local_bb2_shr16_i1654_consumed_1_NO_SHIFT_REG | ~(local_bb2_shr16_i1654_stall_in_1)) & local_bb2_align_0_i1689_stall_local);
		local_bb2_lnot23_i1661_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1689_inputs_ready & (local_bb2_lnot23_i1661_consumed_0_NO_SHIFT_REG | ~(local_bb2_lnot23_i1661_stall_in)) & local_bb2_align_0_i1689_stall_local);
		local_bb2_cmp27_i1663_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1689_inputs_ready & (local_bb2_cmp27_i1663_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp27_i1663_stall_in)) & local_bb2_align_0_i1689_stall_local);
		local_bb2_align_0_i1689_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1689_inputs_ready & (local_bb2_align_0_i1689_consumed_0_NO_SHIFT_REG | ~(local_bb2_align_0_i1689_stall_in)) & local_bb2_align_0_i1689_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_and35_i1664_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1664_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and35_i1664_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1664_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and35_i1664_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1664_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1664_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1664_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_and35_i1664_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_and35_i1664_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_and35_i1664_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_and35_i1664_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_and35_i1664_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2_and35_i1664_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2_and35_i1664_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_and35_i1664_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_and35_i1664_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_and35_i1664_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_and35_i1664_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_and35_i1664_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and35_i1664_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and35_i1664_0_NO_SHIFT_REG = rnode_175to176_bb2_and35_i1664_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_and35_i1664_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and35_i1664_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shl65_i1135_stall_local;
wire [31:0] local_bb2_shl65_i1135;

assign local_bb2_shl65_i1135 = (local_bb2_or64_i1134 | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp69_i1139_stall_local;
wire local_bb2_cmp69_i1139;

assign local_bb2_cmp69_i1139 = (local_bb2_and68_i1138 > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_not_i1123_stall_local;
wire local_bb2_lnot30_not_i1123;

assign local_bb2_lnot30_not_i1123 = (local_bb2_lnot30_i1119 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i1132_stall_local;
wire [31:0] local_bb2_shl_i1132;

assign local_bb2_shl_i1132 = (local_bb2_or_i1131 | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and35_i1115_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1115_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and35_i1115_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1115_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and35_i1115_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1115_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1115_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i1115_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and35_i1115_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and35_i1115_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and35_i1115_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and35_i1115_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and35_i1115_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2_and35_i1115_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2_and35_i1115_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and35_i1115_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and35_i1115_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and35_i1115_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and35_i1115_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and35_i1115_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_and35_i1115_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and35_i1115_0_NO_SHIFT_REG = rnode_174to175_bb2_and35_i1115_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and35_i1115_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and35_i1115_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shl65_i123_stall_local;
wire [31:0] local_bb2_shl65_i123;

assign local_bb2_shl65_i123 = (local_bb2_or64_i122 | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp69_i127_stall_local;
wire local_bb2_cmp69_i127;

assign local_bb2_cmp69_i127 = (local_bb2_and68_i126 > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_not_i111_stall_local;
wire local_bb2_lnot30_not_i111;

assign local_bb2_lnot30_not_i111 = (local_bb2_lnot30_i107 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i120_stall_local;
wire [31:0] local_bb2_shl_i120;

assign local_bb2_shl_i120 = (local_bb2_or_i119 | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and35_i103_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i103_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and35_i103_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i103_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and35_i103_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i103_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i103_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and35_i103_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and35_i103_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and35_i103_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and35_i103_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and35_i103_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and35_i103_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2_and35_i103_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2_and35_i103_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and35_i103_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and35_i103_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and35_i103_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and35_i103_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and35_i103_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_and35_i103_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and35_i103_0_NO_SHIFT_REG = rnode_174to175_bb2_and35_i103_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and35_i103_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and35_i103_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i642_valid_out_1;
wire local_bb2_shr16_i642_stall_in_1;
 reg local_bb2_shr16_i642_consumed_1_NO_SHIFT_REG;
wire local_bb2_lnot23_i649_valid_out;
wire local_bb2_lnot23_i649_stall_in;
 reg local_bb2_lnot23_i649_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp27_i651_valid_out;
wire local_bb2_cmp27_i651_stall_in;
 reg local_bb2_cmp27_i651_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i671_valid_out;
wire local_bb2_align_0_i671_stall_in;
 reg local_bb2_align_0_i671_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i671_inputs_ready;
wire local_bb2_align_0_i671_stall_local;
wire [31:0] local_bb2_align_0_i671;

assign local_bb2_align_0_i671_inputs_ready = (rnode_171to172_bb2__22_i640_0_valid_out_0_NO_SHIFT_REG & rnode_171to172_bb2__23_i641_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_align_0_i671 = (local_bb2_cmp70_i ? 32'h1F : local_bb2_and69_i);
assign local_bb2_shr16_i642_valid_out_1 = 1'b1;
assign local_bb2_lnot23_i649_valid_out = 1'b1;
assign local_bb2_cmp27_i651_valid_out = 1'b1;
assign local_bb2_align_0_i671_valid_out = 1'b1;
assign rnode_171to172_bb2__22_i640_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__23_i641_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_shr16_i642_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lnot23_i649_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp27_i651_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_align_0_i671_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_shr16_i642_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i671_inputs_ready & (local_bb2_shr16_i642_consumed_1_NO_SHIFT_REG | ~(local_bb2_shr16_i642_stall_in_1)) & local_bb2_align_0_i671_stall_local);
		local_bb2_lnot23_i649_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i671_inputs_ready & (local_bb2_lnot23_i649_consumed_0_NO_SHIFT_REG | ~(local_bb2_lnot23_i649_stall_in)) & local_bb2_align_0_i671_stall_local);
		local_bb2_cmp27_i651_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i671_inputs_ready & (local_bb2_cmp27_i651_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp27_i651_stall_in)) & local_bb2_align_0_i671_stall_local);
		local_bb2_align_0_i671_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i671_inputs_ready & (local_bb2_align_0_i671_consumed_0_NO_SHIFT_REG | ~(local_bb2_align_0_i671_stall_in)) & local_bb2_align_0_i671_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_and35_i652_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i652_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and35_i652_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i652_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and35_i652_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i652_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i652_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i652_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_and35_i652_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_and35_i652_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_and35_i652_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_and35_i652_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_and35_i652_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2_and35_i652_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2_and35_i652_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_and35_i652_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_and35_i652_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_and35_i652_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_and35_i652_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_and35_i652_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and35_i652_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and35_i652_0_NO_SHIFT_REG = rnode_175to176_bb2_and35_i652_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_and35_i652_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and35_i652_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_shr16_i1654_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1654_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i1654_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1654_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1654_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i1654_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1654_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i1654_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1654_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1654_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1654_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_shr16_i1654_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_shr16_i1654_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_shr16_i1654_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_shr16_i1654_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_shr16_i1654_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_shr16_i1654),
	.data_out(rnode_172to173_bb2_shr16_i1654_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_shr16_i1654_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_shr16_i1654_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2_shr16_i1654_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_shr16_i1654_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_shr16_i1654_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr16_i1654_stall_in_1 = 1'b0;
assign rnode_172to173_bb2_shr16_i1654_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_shr16_i1654_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i1654_0_NO_SHIFT_REG = rnode_172to173_bb2_shr16_i1654_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_shr16_i1654_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i1654_1_NO_SHIFT_REG = rnode_172to173_bb2_shr16_i1654_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_lnot23_i1661_0_valid_out_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1661_0_stall_in_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1661_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1661_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1661_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1661_0_valid_out_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1661_0_stall_in_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1661_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_lnot23_i1661_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_lnot23_i1661_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_lnot23_i1661_0_stall_in_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_lnot23_i1661_0_valid_out_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_lnot23_i1661_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_lnot23_i1661),
	.data_out(rnode_172to173_bb2_lnot23_i1661_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_lnot23_i1661_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_lnot23_i1661_0_reg_173_fifo.DATA_WIDTH = 1;
defparam rnode_172to173_bb2_lnot23_i1661_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_lnot23_i1661_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_lnot23_i1661_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lnot23_i1661_stall_in = 1'b0;
assign rnode_172to173_bb2_lnot23_i1661_0_NO_SHIFT_REG = rnode_172to173_bb2_lnot23_i1661_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_lnot23_i1661_0_stall_in_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_lnot23_i1661_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_cmp27_i1663_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1663_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_cmp27_i1663_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_cmp27_i1663_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_cmp27_i1663_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_cmp27_i1663_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_cmp27_i1663_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_cmp27_i1663),
	.data_out(rnode_172to173_bb2_cmp27_i1663_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_cmp27_i1663_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_cmp27_i1663_0_reg_173_fifo.DATA_WIDTH = 1;
defparam rnode_172to173_bb2_cmp27_i1663_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_cmp27_i1663_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_cmp27_i1663_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp27_i1663_stall_in = 1'b0;
assign rnode_172to173_bb2_cmp27_i1663_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i1663_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i1663_0_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i1663_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_cmp27_i1663_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i1663_1_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i1663_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_cmp27_i1663_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i1663_2_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i1663_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_align_0_i1689_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1689_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1689_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1689_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1689_3_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1689_4_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1689_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1689_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_align_0_i1689_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_align_0_i1689_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_align_0_i1689_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_align_0_i1689_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_align_0_i1689_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_align_0_i1689),
	.data_out(rnode_172to173_bb2_align_0_i1689_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_align_0_i1689_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_align_0_i1689_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2_align_0_i1689_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_align_0_i1689_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_align_0_i1689_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_align_0_i1689_stall_in = 1'b0;
assign rnode_172to173_bb2_align_0_i1689_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1689_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1689_0_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1689_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i1689_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1689_1_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1689_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i1689_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1689_2_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1689_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i1689_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1689_3_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1689_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i1689_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1689_4_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1689_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i1105_valid_out_1;
wire local_bb2_shr16_i1105_stall_in_1;
 reg local_bb2_shr16_i1105_consumed_1_NO_SHIFT_REG;
wire local_bb2_lnot23_i1112_valid_out;
wire local_bb2_lnot23_i1112_stall_in;
 reg local_bb2_lnot23_i1112_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp27_i1114_valid_out;
wire local_bb2_cmp27_i1114_stall_in;
 reg local_bb2_cmp27_i1114_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i1140_valid_out;
wire local_bb2_align_0_i1140_stall_in;
 reg local_bb2_align_0_i1140_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i1140_inputs_ready;
wire local_bb2_align_0_i1140_stall_local;
wire [31:0] local_bb2_align_0_i1140;

assign local_bb2_align_0_i1140_inputs_ready = (rnode_171to172_bb2__22_i1103_0_valid_out_0_NO_SHIFT_REG & rnode_171to172_bb2__23_i1104_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_align_0_i1140 = (local_bb2_cmp69_i1139 ? 32'h1F : local_bb2_and68_i1138);
assign local_bb2_shr16_i1105_valid_out_1 = 1'b1;
assign local_bb2_lnot23_i1112_valid_out = 1'b1;
assign local_bb2_cmp27_i1114_valid_out = 1'b1;
assign local_bb2_align_0_i1140_valid_out = 1'b1;
assign rnode_171to172_bb2__22_i1103_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__23_i1104_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_shr16_i1105_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lnot23_i1112_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp27_i1114_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_align_0_i1140_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_shr16_i1105_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i1140_inputs_ready & (local_bb2_shr16_i1105_consumed_1_NO_SHIFT_REG | ~(local_bb2_shr16_i1105_stall_in_1)) & local_bb2_align_0_i1140_stall_local);
		local_bb2_lnot23_i1112_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1140_inputs_ready & (local_bb2_lnot23_i1112_consumed_0_NO_SHIFT_REG | ~(local_bb2_lnot23_i1112_stall_in)) & local_bb2_align_0_i1140_stall_local);
		local_bb2_cmp27_i1114_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1140_inputs_ready & (local_bb2_cmp27_i1114_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp27_i1114_stall_in)) & local_bb2_align_0_i1140_stall_local);
		local_bb2_align_0_i1140_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1140_inputs_ready & (local_bb2_align_0_i1140_consumed_0_NO_SHIFT_REG | ~(local_bb2_align_0_i1140_stall_in)) & local_bb2_align_0_i1140_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_and35_i1115_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1115_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and35_i1115_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1115_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and35_i1115_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1115_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1115_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i1115_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_and35_i1115_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_and35_i1115_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_and35_i1115_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_and35_i1115_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_and35_i1115_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2_and35_i1115_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2_and35_i1115_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_and35_i1115_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_and35_i1115_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_and35_i1115_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_and35_i1115_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_and35_i1115_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and35_i1115_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and35_i1115_0_NO_SHIFT_REG = rnode_175to176_bb2_and35_i1115_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_and35_i1115_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and35_i1115_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i93_valid_out_1;
wire local_bb2_shr16_i93_stall_in_1;
 reg local_bb2_shr16_i93_consumed_1_NO_SHIFT_REG;
wire local_bb2_lnot23_i100_valid_out;
wire local_bb2_lnot23_i100_stall_in;
 reg local_bb2_lnot23_i100_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp27_i102_valid_out;
wire local_bb2_cmp27_i102_stall_in;
 reg local_bb2_cmp27_i102_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i128_valid_out;
wire local_bb2_align_0_i128_stall_in;
 reg local_bb2_align_0_i128_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i128_inputs_ready;
wire local_bb2_align_0_i128_stall_local;
wire [31:0] local_bb2_align_0_i128;

assign local_bb2_align_0_i128_inputs_ready = (rnode_171to172_bb2__22_i91_0_valid_out_0_NO_SHIFT_REG & rnode_171to172_bb2__23_i92_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_align_0_i128 = (local_bb2_cmp69_i127 ? 32'h1F : local_bb2_and68_i126);
assign local_bb2_shr16_i93_valid_out_1 = 1'b1;
assign local_bb2_lnot23_i100_valid_out = 1'b1;
assign local_bb2_cmp27_i102_valid_out = 1'b1;
assign local_bb2_align_0_i128_valid_out = 1'b1;
assign rnode_171to172_bb2__22_i91_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_171to172_bb2__23_i92_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_shr16_i93_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lnot23_i100_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp27_i102_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_align_0_i128_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_shr16_i93_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i128_inputs_ready & (local_bb2_shr16_i93_consumed_1_NO_SHIFT_REG | ~(local_bb2_shr16_i93_stall_in_1)) & local_bb2_align_0_i128_stall_local);
		local_bb2_lnot23_i100_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i128_inputs_ready & (local_bb2_lnot23_i100_consumed_0_NO_SHIFT_REG | ~(local_bb2_lnot23_i100_stall_in)) & local_bb2_align_0_i128_stall_local);
		local_bb2_cmp27_i102_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i128_inputs_ready & (local_bb2_cmp27_i102_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp27_i102_stall_in)) & local_bb2_align_0_i128_stall_local);
		local_bb2_align_0_i128_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i128_inputs_ready & (local_bb2_align_0_i128_consumed_0_NO_SHIFT_REG | ~(local_bb2_align_0_i128_stall_in)) & local_bb2_align_0_i128_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_and35_i103_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i103_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and35_i103_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i103_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and35_i103_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i103_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i103_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and35_i103_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_and35_i103_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_and35_i103_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_and35_i103_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_and35_i103_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_and35_i103_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2_and35_i103_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2_and35_i103_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_and35_i103_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_and35_i103_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_and35_i103_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_and35_i103_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_and35_i103_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and35_i103_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and35_i103_0_NO_SHIFT_REG = rnode_175to176_bb2_and35_i103_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_and35_i103_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and35_i103_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_shr16_i642_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i642_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i642_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i642_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i642_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i642_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i642_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i642_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i642_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i642_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i642_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_shr16_i642_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_shr16_i642_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_shr16_i642_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_shr16_i642_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_shr16_i642_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_shr16_i642),
	.data_out(rnode_172to173_bb2_shr16_i642_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_shr16_i642_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_shr16_i642_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2_shr16_i642_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_shr16_i642_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_shr16_i642_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr16_i642_stall_in_1 = 1'b0;
assign rnode_172to173_bb2_shr16_i642_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_shr16_i642_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i642_0_NO_SHIFT_REG = rnode_172to173_bb2_shr16_i642_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_shr16_i642_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i642_1_NO_SHIFT_REG = rnode_172to173_bb2_shr16_i642_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_lnot23_i649_0_valid_out_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i649_0_stall_in_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i649_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i649_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i649_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i649_0_valid_out_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i649_0_stall_in_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i649_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_lnot23_i649_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_lnot23_i649_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_lnot23_i649_0_stall_in_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_lnot23_i649_0_valid_out_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_lnot23_i649_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_lnot23_i649),
	.data_out(rnode_172to173_bb2_lnot23_i649_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_lnot23_i649_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_lnot23_i649_0_reg_173_fifo.DATA_WIDTH = 1;
defparam rnode_172to173_bb2_lnot23_i649_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_lnot23_i649_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_lnot23_i649_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lnot23_i649_stall_in = 1'b0;
assign rnode_172to173_bb2_lnot23_i649_0_NO_SHIFT_REG = rnode_172to173_bb2_lnot23_i649_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_lnot23_i649_0_stall_in_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_lnot23_i649_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_cmp27_i651_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i651_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_cmp27_i651_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_cmp27_i651_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_cmp27_i651_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_cmp27_i651_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_cmp27_i651_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_cmp27_i651),
	.data_out(rnode_172to173_bb2_cmp27_i651_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_cmp27_i651_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_cmp27_i651_0_reg_173_fifo.DATA_WIDTH = 1;
defparam rnode_172to173_bb2_cmp27_i651_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_cmp27_i651_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_cmp27_i651_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp27_i651_stall_in = 1'b0;
assign rnode_172to173_bb2_cmp27_i651_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i651_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i651_0_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i651_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_cmp27_i651_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i651_1_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i651_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_cmp27_i651_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i651_2_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i651_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_align_0_i671_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i671_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i671_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i671_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i671_3_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i671_4_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i671_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i671_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_align_0_i671_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_align_0_i671_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_align_0_i671_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_align_0_i671_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_align_0_i671_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_align_0_i671),
	.data_out(rnode_172to173_bb2_align_0_i671_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_align_0_i671_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_align_0_i671_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2_align_0_i671_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_align_0_i671_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_align_0_i671_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_align_0_i671_stall_in = 1'b0;
assign rnode_172to173_bb2_align_0_i671_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i671_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i671_0_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i671_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i671_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i671_1_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i671_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i671_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i671_2_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i671_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i671_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i671_3_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i671_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i671_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i671_4_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i671_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and17_i1655_stall_local;
wire [31:0] local_bb2_and17_i1655;

assign local_bb2_and17_i1655 = (rnode_172to173_bb2_shr16_i1654_0_NO_SHIFT_REG & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_shr16_i1654_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1654_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_shr16_i1654_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1654_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_shr16_i1654_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1654_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1654_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1654_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_shr16_i1654_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_shr16_i1654_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_shr16_i1654_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_shr16_i1654_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_shr16_i1654_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_172to173_bb2_shr16_i1654_1_NO_SHIFT_REG),
	.data_out(rnode_173to175_bb2_shr16_i1654_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_shr16_i1654_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_shr16_i1654_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_173to175_bb2_shr16_i1654_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_shr16_i1654_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_shr16_i1654_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i1654_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_shr16_i1654_0_NO_SHIFT_REG = rnode_173to175_bb2_shr16_i1654_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_shr16_i1654_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_shr16_i1654_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2__28_i1685_stall_local;
wire [31:0] local_bb2__28_i1685;

assign local_bb2__28_i1685 = (rnode_172to173_bb2_lnot23_i1661_0_NO_SHIFT_REG ? 32'h0 : local_bb2_shl66_i1684);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_i1671_stall_local;
wire local_bb2_brmerge_not_i1671;

assign local_bb2_brmerge_not_i1671 = (rnode_172to173_bb2_cmp27_i1663_0_NO_SHIFT_REG & local_bb2_lnot33_not_i1670);

// This section implements an unregistered operation.
// 
wire local_bb2_and94_i1697_stall_local;
wire [31:0] local_bb2_and94_i1697;

assign local_bb2_and94_i1697 = (rnode_172to173_bb2_align_0_i1689_0_NO_SHIFT_REG & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb2_and96_i1699_stall_local;
wire [31:0] local_bb2_and96_i1699;

assign local_bb2_and96_i1699 = (rnode_172to173_bb2_align_0_i1689_1_NO_SHIFT_REG & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and116_i1715_stall_local;
wire [31:0] local_bb2_and116_i1715;

assign local_bb2_and116_i1715 = (rnode_172to173_bb2_align_0_i1689_2_NO_SHIFT_REG & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_and131_i1721_stall_local;
wire [31:0] local_bb2_and131_i1721;

assign local_bb2_and131_i1721 = (rnode_172to173_bb2_align_0_i1689_3_NO_SHIFT_REG & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and150_i1726_stall_local;
wire [31:0] local_bb2_and150_i1726;

assign local_bb2_and150_i1726 = (rnode_172to173_bb2_align_0_i1689_4_NO_SHIFT_REG & 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_shr16_i1105_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1105_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i1105_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1105_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1105_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i1105_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1105_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i1105_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1105_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1105_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i1105_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_shr16_i1105_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_shr16_i1105_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_shr16_i1105_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_shr16_i1105_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_shr16_i1105_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_shr16_i1105),
	.data_out(rnode_172to173_bb2_shr16_i1105_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_shr16_i1105_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_shr16_i1105_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2_shr16_i1105_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_shr16_i1105_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_shr16_i1105_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr16_i1105_stall_in_1 = 1'b0;
assign rnode_172to173_bb2_shr16_i1105_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_shr16_i1105_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i1105_0_NO_SHIFT_REG = rnode_172to173_bb2_shr16_i1105_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_shr16_i1105_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i1105_1_NO_SHIFT_REG = rnode_172to173_bb2_shr16_i1105_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_lnot23_i1112_0_valid_out_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1112_0_stall_in_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1112_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1112_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1112_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1112_0_valid_out_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1112_0_stall_in_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i1112_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_lnot23_i1112_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_lnot23_i1112_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_lnot23_i1112_0_stall_in_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_lnot23_i1112_0_valid_out_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_lnot23_i1112_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_lnot23_i1112),
	.data_out(rnode_172to173_bb2_lnot23_i1112_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_lnot23_i1112_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_lnot23_i1112_0_reg_173_fifo.DATA_WIDTH = 1;
defparam rnode_172to173_bb2_lnot23_i1112_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_lnot23_i1112_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_lnot23_i1112_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lnot23_i1112_stall_in = 1'b0;
assign rnode_172to173_bb2_lnot23_i1112_0_NO_SHIFT_REG = rnode_172to173_bb2_lnot23_i1112_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_lnot23_i1112_0_stall_in_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_lnot23_i1112_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_cmp27_i1114_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i1114_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_cmp27_i1114_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_cmp27_i1114_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_cmp27_i1114_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_cmp27_i1114_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_cmp27_i1114_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_cmp27_i1114),
	.data_out(rnode_172to173_bb2_cmp27_i1114_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_cmp27_i1114_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_cmp27_i1114_0_reg_173_fifo.DATA_WIDTH = 1;
defparam rnode_172to173_bb2_cmp27_i1114_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_cmp27_i1114_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_cmp27_i1114_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp27_i1114_stall_in = 1'b0;
assign rnode_172to173_bb2_cmp27_i1114_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i1114_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i1114_0_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i1114_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_cmp27_i1114_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i1114_1_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i1114_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_cmp27_i1114_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i1114_2_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i1114_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_align_0_i1140_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1140_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1140_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1140_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1140_3_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1140_4_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i1140_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i1140_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_align_0_i1140_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_align_0_i1140_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_align_0_i1140_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_align_0_i1140_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_align_0_i1140_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_align_0_i1140),
	.data_out(rnode_172to173_bb2_align_0_i1140_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_align_0_i1140_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_align_0_i1140_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2_align_0_i1140_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_align_0_i1140_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_align_0_i1140_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_align_0_i1140_stall_in = 1'b0;
assign rnode_172to173_bb2_align_0_i1140_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1140_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1140_0_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1140_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i1140_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1140_1_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1140_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i1140_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1140_2_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1140_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i1140_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1140_3_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1140_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i1140_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i1140_4_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i1140_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_shr16_i93_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i93_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i93_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i93_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i93_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i93_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i93_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_shr16_i93_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i93_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i93_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_shr16_i93_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_shr16_i93_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_shr16_i93_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_shr16_i93_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_shr16_i93_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_shr16_i93_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_shr16_i93),
	.data_out(rnode_172to173_bb2_shr16_i93_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_shr16_i93_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_shr16_i93_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2_shr16_i93_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_shr16_i93_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_shr16_i93_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr16_i93_stall_in_1 = 1'b0;
assign rnode_172to173_bb2_shr16_i93_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_shr16_i93_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i93_0_NO_SHIFT_REG = rnode_172to173_bb2_shr16_i93_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_shr16_i93_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i93_1_NO_SHIFT_REG = rnode_172to173_bb2_shr16_i93_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_lnot23_i100_0_valid_out_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i100_0_stall_in_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i100_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i100_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i100_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i100_0_valid_out_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i100_0_stall_in_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_lnot23_i100_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_lnot23_i100_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_lnot23_i100_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_lnot23_i100_0_stall_in_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_lnot23_i100_0_valid_out_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_lnot23_i100_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_lnot23_i100),
	.data_out(rnode_172to173_bb2_lnot23_i100_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_lnot23_i100_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_lnot23_i100_0_reg_173_fifo.DATA_WIDTH = 1;
defparam rnode_172to173_bb2_lnot23_i100_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_lnot23_i100_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_lnot23_i100_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lnot23_i100_stall_in = 1'b0;
assign rnode_172to173_bb2_lnot23_i100_0_NO_SHIFT_REG = rnode_172to173_bb2_lnot23_i100_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_lnot23_i100_0_stall_in_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_lnot23_i100_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_cmp27_i102_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_cmp27_i102_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_cmp27_i102_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_cmp27_i102_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_cmp27_i102_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_cmp27_i102_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_cmp27_i102_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_cmp27_i102),
	.data_out(rnode_172to173_bb2_cmp27_i102_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_cmp27_i102_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_cmp27_i102_0_reg_173_fifo.DATA_WIDTH = 1;
defparam rnode_172to173_bb2_cmp27_i102_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_cmp27_i102_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_cmp27_i102_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp27_i102_stall_in = 1'b0;
assign rnode_172to173_bb2_cmp27_i102_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i102_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i102_0_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i102_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_cmp27_i102_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i102_1_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i102_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_cmp27_i102_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_cmp27_i102_2_NO_SHIFT_REG = rnode_172to173_bb2_cmp27_i102_0_reg_173_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_172to173_bb2_align_0_i128_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i128_0_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i128_1_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i128_2_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i128_3_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i128_4_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_reg_173_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_172to173_bb2_align_0_i128_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_valid_out_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_stall_in_0_reg_173_NO_SHIFT_REG;
 logic rnode_172to173_bb2_align_0_i128_0_stall_out_reg_173_NO_SHIFT_REG;

acl_data_fifo rnode_172to173_bb2_align_0_i128_0_reg_173_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_172to173_bb2_align_0_i128_0_reg_173_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_172to173_bb2_align_0_i128_0_stall_in_0_reg_173_NO_SHIFT_REG),
	.valid_out(rnode_172to173_bb2_align_0_i128_0_valid_out_0_reg_173_NO_SHIFT_REG),
	.stall_out(rnode_172to173_bb2_align_0_i128_0_stall_out_reg_173_NO_SHIFT_REG),
	.data_in(local_bb2_align_0_i128),
	.data_out(rnode_172to173_bb2_align_0_i128_0_reg_173_NO_SHIFT_REG)
);

defparam rnode_172to173_bb2_align_0_i128_0_reg_173_fifo.DEPTH = 1;
defparam rnode_172to173_bb2_align_0_i128_0_reg_173_fifo.DATA_WIDTH = 32;
defparam rnode_172to173_bb2_align_0_i128_0_reg_173_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_172to173_bb2_align_0_i128_0_reg_173_fifo.IMPL = "shift_reg";

assign rnode_172to173_bb2_align_0_i128_0_reg_173_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_align_0_i128_stall_in = 1'b0;
assign rnode_172to173_bb2_align_0_i128_0_stall_in_0_reg_173_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i128_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i128_0_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i128_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i128_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i128_1_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i128_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i128_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i128_2_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i128_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i128_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i128_3_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i128_0_reg_173_NO_SHIFT_REG;
assign rnode_172to173_bb2_align_0_i128_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_align_0_i128_4_NO_SHIFT_REG = rnode_172to173_bb2_align_0_i128_0_reg_173_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and17_i643_stall_local;
wire [31:0] local_bb2_and17_i643;

assign local_bb2_and17_i643 = (rnode_172to173_bb2_shr16_i642_0_NO_SHIFT_REG & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_shr16_i642_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i642_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_shr16_i642_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i642_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_shr16_i642_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i642_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i642_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i642_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_shr16_i642_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_shr16_i642_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_shr16_i642_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_shr16_i642_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_shr16_i642_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_172to173_bb2_shr16_i642_1_NO_SHIFT_REG),
	.data_out(rnode_173to175_bb2_shr16_i642_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_shr16_i642_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_shr16_i642_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_173to175_bb2_shr16_i642_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_shr16_i642_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_shr16_i642_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i642_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_shr16_i642_0_NO_SHIFT_REG = rnode_173to175_bb2_shr16_i642_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_shr16_i642_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_shr16_i642_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2__28_i669_stall_local;
wire [31:0] local_bb2__28_i669;

assign local_bb2__28_i669 = (rnode_172to173_bb2_lnot23_i649_0_NO_SHIFT_REG ? 32'h0 : local_bb2_shl66_i);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_i657_stall_local;
wire local_bb2_brmerge_not_i657;

assign local_bb2_brmerge_not_i657 = (rnode_172to173_bb2_cmp27_i651_0_NO_SHIFT_REG & local_bb2_lnot33_not_i656);

// This section implements an unregistered operation.
// 
wire local_bb2_and94_i_stall_local;
wire [31:0] local_bb2_and94_i;

assign local_bb2_and94_i = (rnode_172to173_bb2_align_0_i671_0_NO_SHIFT_REG & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb2_and96_i_stall_local;
wire [31:0] local_bb2_and96_i;

assign local_bb2_and96_i = (rnode_172to173_bb2_align_0_i671_1_NO_SHIFT_REG & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and116_i_stall_local;
wire [31:0] local_bb2_and116_i;

assign local_bb2_and116_i = (rnode_172to173_bb2_align_0_i671_2_NO_SHIFT_REG & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_and131_i_stall_local;
wire [31:0] local_bb2_and131_i;

assign local_bb2_and131_i = (rnode_172to173_bb2_align_0_i671_3_NO_SHIFT_REG & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and150_i_stall_local;
wire [31:0] local_bb2_and150_i;

assign local_bb2_and150_i = (rnode_172to173_bb2_align_0_i671_4_NO_SHIFT_REG & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i1660_stall_local;
wire local_bb2_lnot_i1660;

assign local_bb2_lnot_i1660 = (local_bb2_and17_i1655 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_i1662_stall_local;
wire local_bb2_cmp25_i1662;

assign local_bb2_cmp25_i1662 = (local_bb2_and17_i1655 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and73_i1690_stall_local;
wire [31:0] local_bb2_and73_i1690;

assign local_bb2_and73_i1690 = (local_bb2__28_i1685 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and76_i1693_stall_local;
wire [31:0] local_bb2_and76_i1693;

assign local_bb2_and76_i1693 = (local_bb2__28_i1685 & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb2_and79_i1695_stall_local;
wire [31:0] local_bb2_and79_i1695;

assign local_bb2_and79_i1695 = (local_bb2__28_i1685 & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and91_i1701_stall_local;
wire [31:0] local_bb2_and91_i1701;

assign local_bb2_and91_i1701 = (local_bb2__28_i1685 & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i1702_stall_local;
wire [31:0] local_bb2_and88_i1702;

assign local_bb2_and88_i1702 = (local_bb2__28_i1685 & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb2_and85_i1703_stall_local;
wire [31:0] local_bb2_and85_i1703;

assign local_bb2_and85_i1703 = (local_bb2__28_i1685 & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u100_stall_local;
wire [31:0] local_bb2_var__u100;

assign local_bb2_var__u100 = (local_bb2__28_i1685 & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_not_i1675_stall_local;
wire local_bb2_brmerge_not_not_i1675;

assign local_bb2_brmerge_not_not_i1675 = (local_bb2_brmerge_not_i1671 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr95_i1698_stall_local;
wire [31:0] local_bb2_shr95_i1698;

assign local_bb2_shr95_i1698 = (local_bb2__28_i1685 >> local_bb2_and94_i1697);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp97_i1700_stall_local;
wire local_bb2_cmp97_i1700;

assign local_bb2_cmp97_i1700 = (local_bb2_and96_i1699 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp117_i1716_stall_local;
wire local_bb2_cmp117_i1716;

assign local_bb2_cmp117_i1716 = (local_bb2_and116_i1715 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp132_not_i1723_stall_local;
wire local_bb2_cmp132_not_i1723;

assign local_bb2_cmp132_not_i1723 = (local_bb2_and131_i1721 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_Pivot20_i1728_stall_local;
wire local_bb2_Pivot20_i1728;

assign local_bb2_Pivot20_i1728 = (local_bb2_and150_i1726 < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_SwitchLeaf_i1729_stall_local;
wire local_bb2_SwitchLeaf_i1729;

assign local_bb2_SwitchLeaf_i1729 = (local_bb2_and150_i1726 == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and17_i1106_stall_local;
wire [31:0] local_bb2_and17_i1106;

assign local_bb2_and17_i1106 = (rnode_172to173_bb2_shr16_i1105_0_NO_SHIFT_REG & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_shr16_i1105_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1105_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_shr16_i1105_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1105_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_shr16_i1105_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1105_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1105_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i1105_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_shr16_i1105_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_shr16_i1105_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_shr16_i1105_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_shr16_i1105_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_shr16_i1105_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_172to173_bb2_shr16_i1105_1_NO_SHIFT_REG),
	.data_out(rnode_173to175_bb2_shr16_i1105_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_shr16_i1105_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_shr16_i1105_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_173to175_bb2_shr16_i1105_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_shr16_i1105_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_shr16_i1105_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i1105_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_shr16_i1105_0_NO_SHIFT_REG = rnode_173to175_bb2_shr16_i1105_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_shr16_i1105_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_shr16_i1105_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2__28_i1136_stall_local;
wire [31:0] local_bb2__28_i1136;

assign local_bb2__28_i1136 = (rnode_172to173_bb2_lnot23_i1112_0_NO_SHIFT_REG ? 32'h0 : local_bb2_shl65_i1135);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_i1122_stall_local;
wire local_bb2_brmerge_not_i1122;

assign local_bb2_brmerge_not_i1122 = (rnode_172to173_bb2_cmp27_i1114_0_NO_SHIFT_REG & local_bb2_lnot33_not_i1121);

// This section implements an unregistered operation.
// 
wire local_bb2_and93_i1148_stall_local;
wire [31:0] local_bb2_and93_i1148;

assign local_bb2_and93_i1148 = (rnode_172to173_bb2_align_0_i1140_0_NO_SHIFT_REG & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb2_and95_i1150_stall_local;
wire [31:0] local_bb2_and95_i1150;

assign local_bb2_and95_i1150 = (rnode_172to173_bb2_align_0_i1140_1_NO_SHIFT_REG & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and115_i1166_stall_local;
wire [31:0] local_bb2_and115_i1166;

assign local_bb2_and115_i1166 = (rnode_172to173_bb2_align_0_i1140_2_NO_SHIFT_REG & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_and130_i1172_stall_local;
wire [31:0] local_bb2_and130_i1172;

assign local_bb2_and130_i1172 = (rnode_172to173_bb2_align_0_i1140_3_NO_SHIFT_REG & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and149_i1177_stall_local;
wire [31:0] local_bb2_and149_i1177;

assign local_bb2_and149_i1177 = (rnode_172to173_bb2_align_0_i1140_4_NO_SHIFT_REG & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and17_i94_stall_local;
wire [31:0] local_bb2_and17_i94;

assign local_bb2_and17_i94 = (rnode_172to173_bb2_shr16_i93_0_NO_SHIFT_REG & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_shr16_i93_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i93_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_shr16_i93_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i93_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_shr16_i93_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i93_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i93_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_shr16_i93_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_shr16_i93_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_shr16_i93_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_shr16_i93_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_shr16_i93_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_shr16_i93_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_172to173_bb2_shr16_i93_1_NO_SHIFT_REG),
	.data_out(rnode_173to175_bb2_shr16_i93_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_shr16_i93_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_shr16_i93_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_173to175_bb2_shr16_i93_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_shr16_i93_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_shr16_i93_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_172to173_bb2_shr16_i93_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_shr16_i93_0_NO_SHIFT_REG = rnode_173to175_bb2_shr16_i93_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_shr16_i93_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_shr16_i93_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2__28_i124_stall_local;
wire [31:0] local_bb2__28_i124;

assign local_bb2__28_i124 = (rnode_172to173_bb2_lnot23_i100_0_NO_SHIFT_REG ? 32'h0 : local_bb2_shl65_i123);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_i110_stall_local;
wire local_bb2_brmerge_not_i110;

assign local_bb2_brmerge_not_i110 = (rnode_172to173_bb2_cmp27_i102_0_NO_SHIFT_REG & local_bb2_lnot33_not_i109);

// This section implements an unregistered operation.
// 
wire local_bb2_and93_i136_stall_local;
wire [31:0] local_bb2_and93_i136;

assign local_bb2_and93_i136 = (rnode_172to173_bb2_align_0_i128_0_NO_SHIFT_REG & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb2_and95_i138_stall_local;
wire [31:0] local_bb2_and95_i138;

assign local_bb2_and95_i138 = (rnode_172to173_bb2_align_0_i128_1_NO_SHIFT_REG & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and115_i154_stall_local;
wire [31:0] local_bb2_and115_i154;

assign local_bb2_and115_i154 = (rnode_172to173_bb2_align_0_i128_2_NO_SHIFT_REG & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_and130_i160_stall_local;
wire [31:0] local_bb2_and130_i160;

assign local_bb2_and130_i160 = (rnode_172to173_bb2_align_0_i128_3_NO_SHIFT_REG & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and149_i165_stall_local;
wire [31:0] local_bb2_and149_i165;

assign local_bb2_and149_i165 = (rnode_172to173_bb2_align_0_i128_4_NO_SHIFT_REG & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i648_stall_local;
wire local_bb2_lnot_i648;

assign local_bb2_lnot_i648 = (local_bb2_and17_i643 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_i650_stall_local;
wire local_bb2_cmp25_i650;

assign local_bb2_cmp25_i650 = (local_bb2_and17_i643 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and73_i_stall_local;
wire [31:0] local_bb2_and73_i;

assign local_bb2_and73_i = (local_bb2__28_i669 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and76_i_stall_local;
wire [31:0] local_bb2_and76_i;

assign local_bb2_and76_i = (local_bb2__28_i669 & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb2_and79_i_stall_local;
wire [31:0] local_bb2_and79_i;

assign local_bb2_and79_i = (local_bb2__28_i669 & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and91_i_stall_local;
wire [31:0] local_bb2_and91_i;

assign local_bb2_and91_i = (local_bb2__28_i669 & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and88_i673_stall_local;
wire [31:0] local_bb2_and88_i673;

assign local_bb2_and88_i673 = (local_bb2__28_i669 & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb2_and85_i_stall_local;
wire [31:0] local_bb2_and85_i;

assign local_bb2_and85_i = (local_bb2__28_i669 & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u101_stall_local;
wire [31:0] local_bb2_var__u101;

assign local_bb2_var__u101 = (local_bb2__28_i669 & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_not_i661_stall_local;
wire local_bb2_brmerge_not_not_i661;

assign local_bb2_brmerge_not_not_i661 = (local_bb2_brmerge_not_i657 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr95_i_stall_local;
wire [31:0] local_bb2_shr95_i;

assign local_bb2_shr95_i = (local_bb2__28_i669 >> local_bb2_and94_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp97_i_stall_local;
wire local_bb2_cmp97_i;

assign local_bb2_cmp97_i = (local_bb2_and96_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp117_i_stall_local;
wire local_bb2_cmp117_i;

assign local_bb2_cmp117_i = (local_bb2_and116_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp132_not_i_stall_local;
wire local_bb2_cmp132_not_i;

assign local_bb2_cmp132_not_i = (local_bb2_and131_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_Pivot20_i682_stall_local;
wire local_bb2_Pivot20_i682;

assign local_bb2_Pivot20_i682 = (local_bb2_and150_i < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_SwitchLeaf_i683_stall_local;
wire local_bb2_SwitchLeaf_i683;

assign local_bb2_SwitchLeaf_i683 = (local_bb2_and150_i == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i1682_stall_local;
wire [31:0] local_bb2__27_i1682;

assign local_bb2__27_i1682 = (local_bb2_lnot_i1660 ? 32'h0 : local_bb2_shl_i1681);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_not_i1667_stall_local;
wire local_bb2_cmp25_not_i1667;

assign local_bb2_cmp25_not_i1667 = (local_bb2_cmp25_i1662 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_not_i1673_stall_local;
wire local_bb2_or_cond_not_i1673;

assign local_bb2_or_cond_not_i1673 = (local_bb2_cmp25_i1662 & local_bb2_lnot30_not_i1672);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u102_stall_local;
wire local_bb2_var__u102;

assign local_bb2_var__u102 = (local_bb2_cmp25_i1662 | rnode_172to173_bb2_cmp27_i1663_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and73_tr_i1691_stall_local;
wire [7:0] local_bb2_and73_tr_i1691;

assign local_bb2_and73_tr_i1691 = local_bb2_and73_i1690[7:0];

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i1694_stall_local;
wire local_bb2_cmp77_i1694;

assign local_bb2_cmp77_i1694 = (local_bb2_and76_i1693 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp80_i1696_stall_local;
wire local_bb2_cmp80_i1696;

assign local_bb2_cmp80_i1696 = (local_bb2_and79_i1695 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp92_i1704_stall_local;
wire local_bb2_cmp92_i1704;

assign local_bb2_cmp92_i1704 = (local_bb2_and91_i1701 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp89_i1705_stall_local;
wire local_bb2_cmp89_i1705;

assign local_bb2_cmp89_i1705 = (local_bb2_and88_i1702 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp86_i1706_stall_local;
wire local_bb2_cmp86_i1706;

assign local_bb2_cmp86_i1706 = (local_bb2_and85_i1703 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u103_stall_local;
wire local_bb2_var__u103;

assign local_bb2_var__u103 = (local_bb2_var__u100 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_7_i1676_stall_local;
wire local_bb2_reduction_7_i1676;

assign local_bb2_reduction_7_i1676 = (local_bb2_cmp25_i1662 & local_bb2_brmerge_not_not_i1675);

// This section implements an unregistered operation.
// 
wire local_bb2_and143_i1725_stall_local;
wire [31:0] local_bb2_and143_i1725;

assign local_bb2_and143_i1725 = (local_bb2_shr95_i1698 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr151_i1727_stall_local;
wire [31:0] local_bb2_shr151_i1727;

assign local_bb2_shr151_i1727 = (local_bb2_shr95_i1698 >> local_bb2_and150_i1726);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u104_stall_local;
wire [31:0] local_bb2_var__u104;

assign local_bb2_var__u104 = (local_bb2_shr95_i1698 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and147_i1730_stall_local;
wire [31:0] local_bb2_and147_i1730;

assign local_bb2_and147_i1730 = (local_bb2_shr95_i1698 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i1111_stall_local;
wire local_bb2_lnot_i1111;

assign local_bb2_lnot_i1111 = (local_bb2_and17_i1106 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_i1113_stall_local;
wire local_bb2_cmp25_i1113;

assign local_bb2_cmp25_i1113 = (local_bb2_and17_i1106 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_i1141_stall_local;
wire [31:0] local_bb2_and72_i1141;

assign local_bb2_and72_i1141 = (local_bb2__28_i1136 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i1144_stall_local;
wire [31:0] local_bb2_and75_i1144;

assign local_bb2_and75_i1144 = (local_bb2__28_i1136 & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb2_and78_i1146_stall_local;
wire [31:0] local_bb2_and78_i1146;

assign local_bb2_and78_i1146 = (local_bb2__28_i1136 & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i1152_stall_local;
wire [31:0] local_bb2_and90_i1152;

assign local_bb2_and90_i1152 = (local_bb2__28_i1136 & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and87_i1153_stall_local;
wire [31:0] local_bb2_and87_i1153;

assign local_bb2_and87_i1153 = (local_bb2__28_i1136 & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb2_and84_i1154_stall_local;
wire [31:0] local_bb2_and84_i1154;

assign local_bb2_and84_i1154 = (local_bb2__28_i1136 & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u105_stall_local;
wire [31:0] local_bb2_var__u105;

assign local_bb2_var__u105 = (local_bb2__28_i1136 & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_not_i1126_stall_local;
wire local_bb2_brmerge_not_not_i1126;

assign local_bb2_brmerge_not_not_i1126 = (local_bb2_brmerge_not_i1122 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr94_i1149_stall_local;
wire [31:0] local_bb2_shr94_i1149;

assign local_bb2_shr94_i1149 = (local_bb2__28_i1136 >> local_bb2_and93_i1148);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp96_i1151_stall_local;
wire local_bb2_cmp96_i1151;

assign local_bb2_cmp96_i1151 = (local_bb2_and95_i1150 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp116_i1167_stall_local;
wire local_bb2_cmp116_i1167;

assign local_bb2_cmp116_i1167 = (local_bb2_and115_i1166 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp131_not_i1174_stall_local;
wire local_bb2_cmp131_not_i1174;

assign local_bb2_cmp131_not_i1174 = (local_bb2_and130_i1172 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_Pivot20_i1179_stall_local;
wire local_bb2_Pivot20_i1179;

assign local_bb2_Pivot20_i1179 = (local_bb2_and149_i1177 < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_SwitchLeaf_i1180_stall_local;
wire local_bb2_SwitchLeaf_i1180;

assign local_bb2_SwitchLeaf_i1180 = (local_bb2_and149_i1177 == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i99_stall_local;
wire local_bb2_lnot_i99;

assign local_bb2_lnot_i99 = (local_bb2_and17_i94 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_i101_stall_local;
wire local_bb2_cmp25_i101;

assign local_bb2_cmp25_i101 = (local_bb2_and17_i94 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_i129_stall_local;
wire [31:0] local_bb2_and72_i129;

assign local_bb2_and72_i129 = (local_bb2__28_i124 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i132_stall_local;
wire [31:0] local_bb2_and75_i132;

assign local_bb2_and75_i132 = (local_bb2__28_i124 & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb2_and78_i134_stall_local;
wire [31:0] local_bb2_and78_i134;

assign local_bb2_and78_i134 = (local_bb2__28_i124 & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i140_stall_local;
wire [31:0] local_bb2_and90_i140;

assign local_bb2_and90_i140 = (local_bb2__28_i124 & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and87_i141_stall_local;
wire [31:0] local_bb2_and87_i141;

assign local_bb2_and87_i141 = (local_bb2__28_i124 & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb2_and84_i142_stall_local;
wire [31:0] local_bb2_and84_i142;

assign local_bb2_and84_i142 = (local_bb2__28_i124 & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u106_stall_local;
wire [31:0] local_bb2_var__u106;

assign local_bb2_var__u106 = (local_bb2__28_i124 & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_not_i114_stall_local;
wire local_bb2_brmerge_not_not_i114;

assign local_bb2_brmerge_not_not_i114 = (local_bb2_brmerge_not_i110 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr94_i137_stall_local;
wire [31:0] local_bb2_shr94_i137;

assign local_bb2_shr94_i137 = (local_bb2__28_i124 >> local_bb2_and93_i136);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp96_i139_stall_local;
wire local_bb2_cmp96_i139;

assign local_bb2_cmp96_i139 = (local_bb2_and95_i138 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp116_i155_stall_local;
wire local_bb2_cmp116_i155;

assign local_bb2_cmp116_i155 = (local_bb2_and115_i154 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp131_not_i162_stall_local;
wire local_bb2_cmp131_not_i162;

assign local_bb2_cmp131_not_i162 = (local_bb2_and130_i160 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_Pivot20_i167_stall_local;
wire local_bb2_Pivot20_i167;

assign local_bb2_Pivot20_i167 = (local_bb2_and149_i165 < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_SwitchLeaf_i168_stall_local;
wire local_bb2_SwitchLeaf_i168;

assign local_bb2_SwitchLeaf_i168 = (local_bb2_and149_i165 == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i668_stall_local;
wire [31:0] local_bb2__27_i668;

assign local_bb2__27_i668 = (local_bb2_lnot_i648 ? 32'h0 : local_bb2_shl_i667);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_not_i653_stall_local;
wire local_bb2_cmp25_not_i653;

assign local_bb2_cmp25_not_i653 = (local_bb2_cmp25_i650 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_not_i659_stall_local;
wire local_bb2_or_cond_not_i659;

assign local_bb2_or_cond_not_i659 = (local_bb2_cmp25_i650 & local_bb2_lnot30_not_i658);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u107_stall_local;
wire local_bb2_var__u107;

assign local_bb2_var__u107 = (local_bb2_cmp25_i650 | rnode_172to173_bb2_cmp27_i651_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and73_tr_i_stall_local;
wire [7:0] local_bb2_and73_tr_i;

assign local_bb2_and73_tr_i = local_bb2_and73_i[7:0];

// This section implements an unregistered operation.
// 
wire local_bb2_cmp77_i672_stall_local;
wire local_bb2_cmp77_i672;

assign local_bb2_cmp77_i672 = (local_bb2_and76_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp80_i_stall_local;
wire local_bb2_cmp80_i;

assign local_bb2_cmp80_i = (local_bb2_and79_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp92_i_stall_local;
wire local_bb2_cmp92_i;

assign local_bb2_cmp92_i = (local_bb2_and91_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp89_i_stall_local;
wire local_bb2_cmp89_i;

assign local_bb2_cmp89_i = (local_bb2_and88_i673 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp86_i_stall_local;
wire local_bb2_cmp86_i;

assign local_bb2_cmp86_i = (local_bb2_and85_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u108_stall_local;
wire local_bb2_var__u108;

assign local_bb2_var__u108 = (local_bb2_var__u101 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_7_i662_stall_local;
wire local_bb2_reduction_7_i662;

assign local_bb2_reduction_7_i662 = (local_bb2_cmp25_i650 & local_bb2_brmerge_not_not_i661);

// This section implements an unregistered operation.
// 
wire local_bb2_and143_i_stall_local;
wire [31:0] local_bb2_and143_i;

assign local_bb2_and143_i = (local_bb2_shr95_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr151_i_stall_local;
wire [31:0] local_bb2_shr151_i;

assign local_bb2_shr151_i = (local_bb2_shr95_i >> local_bb2_and150_i);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u109_stall_local;
wire [31:0] local_bb2_var__u109;

assign local_bb2_var__u109 = (local_bb2_shr95_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and147_i_stall_local;
wire [31:0] local_bb2_and147_i;

assign local_bb2_and147_i = (local_bb2_shr95_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i1742_stall_local;
wire [31:0] local_bb2_add_i1742;

assign local_bb2_add_i1742 = (local_bb2__27_i1682 | local_bb2_and37_lobit_i1741);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_i1669_stall_local;
wire local_bb2_or_cond_i1669;

assign local_bb2_or_cond_i1669 = (local_bb2_lnot30_i1668 | local_bb2_cmp25_not_i1667);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i1674_stall_local;
wire local_bb2__24_i1674;

assign local_bb2__24_i1674 = (local_bb2_or_cond_not_i1673 | local_bb2_brmerge_not_i1671);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool75_i1692_stall_local;
wire [7:0] local_bb2_frombool75_i1692;

assign local_bb2_frombool75_i1692 = (local_bb2_and73_tr_i1691 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_v_i1712_stall_local;
wire local_bb2__31_v_i1712;

assign local_bb2__31_v_i1712 = (local_bb2_cmp97_i1700 ? local_bb2_cmp80_i1696 : local_bb2_cmp92_i1704);

// This section implements an unregistered operation.
// 
wire local_bb2__30_v_i1710_stall_local;
wire local_bb2__30_v_i1710;

assign local_bb2__30_v_i1710 = (local_bb2_cmp97_i1700 ? local_bb2_cmp77_i1694 : local_bb2_cmp89_i1705);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool110_i1708_stall_local;
wire [7:0] local_bb2_frombool110_i1708;

assign local_bb2_frombool110_i1708[7:1] = 7'h0;
assign local_bb2_frombool110_i1708[0] = local_bb2_cmp86_i1706;

// This section implements an unregistered operation.
// 
wire local_bb2_or108_i1707_stall_local;
wire [31:0] local_bb2_or108_i1707;

assign local_bb2_or108_i1707[31:1] = 31'h0;
assign local_bb2_or108_i1707[0] = local_bb2_var__u103;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u110_stall_local;
wire [31:0] local_bb2_var__u110;

assign local_bb2_var__u110 = (local_bb2_and147_i1730 | local_bb2_shr95_i1698);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i1133_stall_local;
wire [31:0] local_bb2__27_i1133;

assign local_bb2__27_i1133 = (local_bb2_lnot_i1111 ? 32'h0 : local_bb2_shl_i1132);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_not_i1118_stall_local;
wire local_bb2_cmp25_not_i1118;

assign local_bb2_cmp25_not_i1118 = (local_bb2_cmp25_i1113 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_not_i1124_stall_local;
wire local_bb2_or_cond_not_i1124;

assign local_bb2_or_cond_not_i1124 = (local_bb2_cmp25_i1113 & local_bb2_lnot30_not_i1123);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u111_stall_local;
wire local_bb2_var__u111;

assign local_bb2_var__u111 = (local_bb2_cmp25_i1113 | rnode_172to173_bb2_cmp27_i1114_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_tr_i1142_stall_local;
wire [7:0] local_bb2_and72_tr_i1142;

assign local_bb2_and72_tr_i1142 = local_bb2_and72_i1141[7:0];

// This section implements an unregistered operation.
// 
wire local_bb2_cmp76_i1145_stall_local;
wire local_bb2_cmp76_i1145;

assign local_bb2_cmp76_i1145 = (local_bb2_and75_i1144 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp79_i1147_stall_local;
wire local_bb2_cmp79_i1147;

assign local_bb2_cmp79_i1147 = (local_bb2_and78_i1146 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i1155_stall_local;
wire local_bb2_cmp91_i1155;

assign local_bb2_cmp91_i1155 = (local_bb2_and90_i1152 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp88_i1156_stall_local;
wire local_bb2_cmp88_i1156;

assign local_bb2_cmp88_i1156 = (local_bb2_and87_i1153 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp85_i1157_stall_local;
wire local_bb2_cmp85_i1157;

assign local_bb2_cmp85_i1157 = (local_bb2_and84_i1154 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u112_stall_local;
wire local_bb2_var__u112;

assign local_bb2_var__u112 = (local_bb2_var__u105 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_7_i1127_stall_local;
wire local_bb2_reduction_7_i1127;

assign local_bb2_reduction_7_i1127 = (local_bb2_cmp25_i1113 & local_bb2_brmerge_not_not_i1126);

// This section implements an unregistered operation.
// 
wire local_bb2_and142_i1176_stall_local;
wire [31:0] local_bb2_and142_i1176;

assign local_bb2_and142_i1176 = (local_bb2_shr94_i1149 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr150_i1178_stall_local;
wire [31:0] local_bb2_shr150_i1178;

assign local_bb2_shr150_i1178 = (local_bb2_shr94_i1149 >> local_bb2_and149_i1177);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u113_stall_local;
wire [31:0] local_bb2_var__u113;

assign local_bb2_var__u113 = (local_bb2_shr94_i1149 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and146_i1181_stall_local;
wire [31:0] local_bb2_and146_i1181;

assign local_bb2_and146_i1181 = (local_bb2_shr94_i1149 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i121_stall_local;
wire [31:0] local_bb2__27_i121;

assign local_bb2__27_i121 = (local_bb2_lnot_i99 ? 32'h0 : local_bb2_shl_i120);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_not_i106_stall_local;
wire local_bb2_cmp25_not_i106;

assign local_bb2_cmp25_not_i106 = (local_bb2_cmp25_i101 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_not_i112_stall_local;
wire local_bb2_or_cond_not_i112;

assign local_bb2_or_cond_not_i112 = (local_bb2_cmp25_i101 & local_bb2_lnot30_not_i111);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u114_stall_local;
wire local_bb2_var__u114;

assign local_bb2_var__u114 = (local_bb2_cmp25_i101 | rnode_172to173_bb2_cmp27_i102_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_tr_i130_stall_local;
wire [7:0] local_bb2_and72_tr_i130;

assign local_bb2_and72_tr_i130 = local_bb2_and72_i129[7:0];

// This section implements an unregistered operation.
// 
wire local_bb2_cmp76_i133_stall_local;
wire local_bb2_cmp76_i133;

assign local_bb2_cmp76_i133 = (local_bb2_and75_i132 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp79_i135_stall_local;
wire local_bb2_cmp79_i135;

assign local_bb2_cmp79_i135 = (local_bb2_and78_i134 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i143_stall_local;
wire local_bb2_cmp91_i143;

assign local_bb2_cmp91_i143 = (local_bb2_and90_i140 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp88_i144_stall_local;
wire local_bb2_cmp88_i144;

assign local_bb2_cmp88_i144 = (local_bb2_and87_i141 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp85_i145_stall_local;
wire local_bb2_cmp85_i145;

assign local_bb2_cmp85_i145 = (local_bb2_and84_i142 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u115_stall_local;
wire local_bb2_var__u115;

assign local_bb2_var__u115 = (local_bb2_var__u106 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_7_i115_stall_local;
wire local_bb2_reduction_7_i115;

assign local_bb2_reduction_7_i115 = (local_bb2_cmp25_i101 & local_bb2_brmerge_not_not_i114);

// This section implements an unregistered operation.
// 
wire local_bb2_and142_i164_stall_local;
wire [31:0] local_bb2_and142_i164;

assign local_bb2_and142_i164 = (local_bb2_shr94_i137 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr150_i166_stall_local;
wire [31:0] local_bb2_shr150_i166;

assign local_bb2_shr150_i166 = (local_bb2_shr94_i137 >> local_bb2_and149_i165);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u116_stall_local;
wire [31:0] local_bb2_var__u116;

assign local_bb2_var__u116 = (local_bb2_shr94_i137 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and146_i169_stall_local;
wire [31:0] local_bb2_and146_i169;

assign local_bb2_and146_i169 = (local_bb2_shr94_i137 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i690_stall_local;
wire [31:0] local_bb2_add_i690;

assign local_bb2_add_i690 = (local_bb2__27_i668 | local_bb2_and37_lobit_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_i655_stall_local;
wire local_bb2_or_cond_i655;

assign local_bb2_or_cond_i655 = (local_bb2_lnot30_i654 | local_bb2_cmp25_not_i653);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i660_stall_local;
wire local_bb2__24_i660;

assign local_bb2__24_i660 = (local_bb2_or_cond_not_i659 | local_bb2_brmerge_not_i657);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool75_i_stall_local;
wire [7:0] local_bb2_frombool75_i;

assign local_bb2_frombool75_i = (local_bb2_and73_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_v_i677_stall_local;
wire local_bb2__31_v_i677;

assign local_bb2__31_v_i677 = (local_bb2_cmp97_i ? local_bb2_cmp80_i : local_bb2_cmp92_i);

// This section implements an unregistered operation.
// 
wire local_bb2__30_v_i675_stall_local;
wire local_bb2__30_v_i675;

assign local_bb2__30_v_i675 = (local_bb2_cmp97_i ? local_bb2_cmp77_i672 : local_bb2_cmp89_i);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool110_i_stall_local;
wire [7:0] local_bb2_frombool110_i;

assign local_bb2_frombool110_i[7:1] = 7'h0;
assign local_bb2_frombool110_i[0] = local_bb2_cmp86_i;

// This section implements an unregistered operation.
// 
wire local_bb2_or108_i_stall_local;
wire [31:0] local_bb2_or108_i;

assign local_bb2_or108_i[31:1] = 31'h0;
assign local_bb2_or108_i[0] = local_bb2_var__u108;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u117_stall_local;
wire [31:0] local_bb2_var__u117;

assign local_bb2_var__u117 = (local_bb2_and147_i | local_bb2_shr95_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_8_i1677_stall_local;
wire local_bb2_reduction_8_i1677;

assign local_bb2_reduction_8_i1677 = (rnode_172to173_bb2_cmp27_i1663_1_NO_SHIFT_REG & local_bb2_or_cond_i1669);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i1713_stall_local;
wire [7:0] local_bb2__31_i1713;

assign local_bb2__31_i1713[7:1] = 7'h0;
assign local_bb2__31_i1713[0] = local_bb2__31_v_i1712;

// This section implements an unregistered operation.
// 
wire local_bb2__30_i1711_stall_local;
wire [7:0] local_bb2__30_i1711;

assign local_bb2__30_i1711[7:1] = 7'h0;
assign local_bb2__30_i1711[0] = local_bb2__30_v_i1710;

// This section implements an unregistered operation.
// 
wire local_bb2__29_i1709_stall_local;
wire [7:0] local_bb2__29_i1709;

assign local_bb2__29_i1709 = (local_bb2_cmp97_i1700 ? local_bb2_frombool75_i1692 : local_bb2_frombool110_i1708);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i1714_stall_local;
wire [31:0] local_bb2__32_i1714;

assign local_bb2__32_i1714 = (local_bb2_cmp97_i1700 ? 32'h0 : local_bb2_or108_i1707);

// This section implements an unregistered operation.
// 
wire local_bb2_or1606_i1731_stall_local;
wire [31:0] local_bb2_or1606_i1731;

assign local_bb2_or1606_i1731 = (local_bb2_var__u110 | local_bb2_and143_i1725);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i1193_stall_local;
wire [31:0] local_bb2_add_i1193;

assign local_bb2_add_i1193 = (local_bb2__27_i1133 | local_bb2_and36_lobit_i1192);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_i1120_stall_local;
wire local_bb2_or_cond_i1120;

assign local_bb2_or_cond_i1120 = (local_bb2_lnot30_i1119 | local_bb2_cmp25_not_i1118);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i1125_stall_local;
wire local_bb2__24_i1125;

assign local_bb2__24_i1125 = (local_bb2_or_cond_not_i1124 | local_bb2_brmerge_not_i1122);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool74_i1143_stall_local;
wire [7:0] local_bb2_frombool74_i1143;

assign local_bb2_frombool74_i1143 = (local_bb2_and72_tr_i1142 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_v_i1163_stall_local;
wire local_bb2__31_v_i1163;

assign local_bb2__31_v_i1163 = (local_bb2_cmp96_i1151 ? local_bb2_cmp79_i1147 : local_bb2_cmp91_i1155);

// This section implements an unregistered operation.
// 
wire local_bb2__30_v_i1161_stall_local;
wire local_bb2__30_v_i1161;

assign local_bb2__30_v_i1161 = (local_bb2_cmp96_i1151 ? local_bb2_cmp76_i1145 : local_bb2_cmp88_i1156);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool109_i1159_stall_local;
wire [7:0] local_bb2_frombool109_i1159;

assign local_bb2_frombool109_i1159[7:1] = 7'h0;
assign local_bb2_frombool109_i1159[0] = local_bb2_cmp85_i1157;

// This section implements an unregistered operation.
// 
wire local_bb2_or107_i1158_stall_local;
wire [31:0] local_bb2_or107_i1158;

assign local_bb2_or107_i1158[31:1] = 31'h0;
assign local_bb2_or107_i1158[0] = local_bb2_var__u112;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u118_stall_local;
wire [31:0] local_bb2_var__u118;

assign local_bb2_var__u118 = (local_bb2_and146_i1181 | local_bb2_shr94_i1149);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i181_stall_local;
wire [31:0] local_bb2_add_i181;

assign local_bb2_add_i181 = (local_bb2__27_i121 | local_bb2_and36_lobit_i180);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_i108_stall_local;
wire local_bb2_or_cond_i108;

assign local_bb2_or_cond_i108 = (local_bb2_lnot30_i107 | local_bb2_cmp25_not_i106);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i113_stall_local;
wire local_bb2__24_i113;

assign local_bb2__24_i113 = (local_bb2_or_cond_not_i112 | local_bb2_brmerge_not_i110);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool74_i131_stall_local;
wire [7:0] local_bb2_frombool74_i131;

assign local_bb2_frombool74_i131 = (local_bb2_and72_tr_i130 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_v_i151_stall_local;
wire local_bb2__31_v_i151;

assign local_bb2__31_v_i151 = (local_bb2_cmp96_i139 ? local_bb2_cmp79_i135 : local_bb2_cmp91_i143);

// This section implements an unregistered operation.
// 
wire local_bb2__30_v_i149_stall_local;
wire local_bb2__30_v_i149;

assign local_bb2__30_v_i149 = (local_bb2_cmp96_i139 ? local_bb2_cmp76_i133 : local_bb2_cmp88_i144);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool109_i147_stall_local;
wire [7:0] local_bb2_frombool109_i147;

assign local_bb2_frombool109_i147[7:1] = 7'h0;
assign local_bb2_frombool109_i147[0] = local_bb2_cmp85_i145;

// This section implements an unregistered operation.
// 
wire local_bb2_or107_i146_stall_local;
wire [31:0] local_bb2_or107_i146;

assign local_bb2_or107_i146[31:1] = 31'h0;
assign local_bb2_or107_i146[0] = local_bb2_var__u115;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u119_stall_local;
wire [31:0] local_bb2_var__u119;

assign local_bb2_var__u119 = (local_bb2_and146_i169 | local_bb2_shr94_i137);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_8_i663_stall_local;
wire local_bb2_reduction_8_i663;

assign local_bb2_reduction_8_i663 = (rnode_172to173_bb2_cmp27_i651_1_NO_SHIFT_REG & local_bb2_or_cond_i655);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i678_stall_local;
wire [7:0] local_bb2__31_i678;

assign local_bb2__31_i678[7:1] = 7'h0;
assign local_bb2__31_i678[0] = local_bb2__31_v_i677;

// This section implements an unregistered operation.
// 
wire local_bb2__30_i676_stall_local;
wire [7:0] local_bb2__30_i676;

assign local_bb2__30_i676[7:1] = 7'h0;
assign local_bb2__30_i676[0] = local_bb2__30_v_i675;

// This section implements an unregistered operation.
// 
wire local_bb2__29_i674_stall_local;
wire [7:0] local_bb2__29_i674;

assign local_bb2__29_i674 = (local_bb2_cmp97_i ? local_bb2_frombool75_i : local_bb2_frombool110_i);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i679_stall_local;
wire [31:0] local_bb2__32_i679;

assign local_bb2__32_i679 = (local_bb2_cmp97_i ? 32'h0 : local_bb2_or108_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or1606_i_stall_local;
wire [31:0] local_bb2_or1606_i;

assign local_bb2_or1606_i = (local_bb2_var__u117 | local_bb2_and143_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_9_i1678_stall_local;
wire local_bb2_reduction_9_i1678;

assign local_bb2_reduction_9_i1678 = (local_bb2_reduction_7_i1676 & local_bb2_reduction_8_i1677);

// This section implements an unregistered operation.
// 
wire local_bb2_or1247_i1717_stall_local;
wire [7:0] local_bb2_or1247_i1717;

assign local_bb2_or1247_i1717 = (local_bb2__30_i1711 | local_bb2__29_i1709);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i1719_stall_local;
wire [7:0] local_bb2__33_i1719;

assign local_bb2__33_i1719 = (local_bb2_cmp117_i1716 ? local_bb2__29_i1709 : local_bb2__31_i1713);

// This section implements an unregistered operation.
// 
wire local_bb2_or163_i1732_stall_local;
wire [31:0] local_bb2_or163_i1732;

assign local_bb2_or163_i1732 = (local_bb2_or1606_i1731 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_8_i1128_stall_local;
wire local_bb2_reduction_8_i1128;

assign local_bb2_reduction_8_i1128 = (rnode_172to173_bb2_cmp27_i1114_1_NO_SHIFT_REG & local_bb2_or_cond_i1120);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i1164_stall_local;
wire [7:0] local_bb2__31_i1164;

assign local_bb2__31_i1164[7:1] = 7'h0;
assign local_bb2__31_i1164[0] = local_bb2__31_v_i1163;

// This section implements an unregistered operation.
// 
wire local_bb2__30_i1162_stall_local;
wire [7:0] local_bb2__30_i1162;

assign local_bb2__30_i1162[7:1] = 7'h0;
assign local_bb2__30_i1162[0] = local_bb2__30_v_i1161;

// This section implements an unregistered operation.
// 
wire local_bb2__29_i1160_stall_local;
wire [7:0] local_bb2__29_i1160;

assign local_bb2__29_i1160 = (local_bb2_cmp96_i1151 ? local_bb2_frombool74_i1143 : local_bb2_frombool109_i1159);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i1165_stall_local;
wire [31:0] local_bb2__32_i1165;

assign local_bb2__32_i1165 = (local_bb2_cmp96_i1151 ? 32'h0 : local_bb2_or107_i1158);

// This section implements an unregistered operation.
// 
wire local_bb2_or1596_i1182_stall_local;
wire [31:0] local_bb2_or1596_i1182;

assign local_bb2_or1596_i1182 = (local_bb2_var__u118 | local_bb2_and142_i1176);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_8_i116_stall_local;
wire local_bb2_reduction_8_i116;

assign local_bb2_reduction_8_i116 = (rnode_172to173_bb2_cmp27_i102_1_NO_SHIFT_REG & local_bb2_or_cond_i108);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i152_stall_local;
wire [7:0] local_bb2__31_i152;

assign local_bb2__31_i152[7:1] = 7'h0;
assign local_bb2__31_i152[0] = local_bb2__31_v_i151;

// This section implements an unregistered operation.
// 
wire local_bb2__30_i150_stall_local;
wire [7:0] local_bb2__30_i150;

assign local_bb2__30_i150[7:1] = 7'h0;
assign local_bb2__30_i150[0] = local_bb2__30_v_i149;

// This section implements an unregistered operation.
// 
wire local_bb2__29_i148_stall_local;
wire [7:0] local_bb2__29_i148;

assign local_bb2__29_i148 = (local_bb2_cmp96_i139 ? local_bb2_frombool74_i131 : local_bb2_frombool109_i147);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i153_stall_local;
wire [31:0] local_bb2__32_i153;

assign local_bb2__32_i153 = (local_bb2_cmp96_i139 ? 32'h0 : local_bb2_or107_i146);

// This section implements an unregistered operation.
// 
wire local_bb2_or1596_i170_stall_local;
wire [31:0] local_bb2_or1596_i170;

assign local_bb2_or1596_i170 = (local_bb2_var__u119 | local_bb2_and142_i164);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_9_i664_stall_local;
wire local_bb2_reduction_9_i664;

assign local_bb2_reduction_9_i664 = (local_bb2_reduction_7_i662 & local_bb2_reduction_8_i663);

// This section implements an unregistered operation.
// 
wire local_bb2_or1247_i_stall_local;
wire [7:0] local_bb2_or1247_i;

assign local_bb2_or1247_i = (local_bb2__30_i676 | local_bb2__29_i674);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i681_stall_local;
wire [7:0] local_bb2__33_i681;

assign local_bb2__33_i681 = (local_bb2_cmp117_i ? local_bb2__29_i674 : local_bb2__31_i678);

// This section implements an unregistered operation.
// 
wire local_bb2_or163_i_stall_local;
wire [31:0] local_bb2_or163_i;

assign local_bb2_or163_i = (local_bb2_or1606_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__26_i1679_stall_local;
wire local_bb2__26_i1679;

assign local_bb2__26_i1679 = (local_bb2_reduction_9_i1678 ? local_bb2_cmp38_i1666 : local_bb2__24_i1674);

// This section implements an unregistered operation.
// 
wire local_bb2_or124_i1718_stall_local;
wire [31:0] local_bb2_or124_i1718;

assign local_bb2_or124_i1718[31:8] = 24'h0;
assign local_bb2_or124_i1718[7:0] = local_bb2_or1247_i1717;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u120_stall_local;
wire [7:0] local_bb2_var__u120;

assign local_bb2_var__u120 = (local_bb2__33_i1719 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__37_v_i1733_stall_local;
wire [31:0] local_bb2__37_v_i1733;

assign local_bb2__37_v_i1733 = (local_bb2_Pivot20_i1728 ? 32'h0 : local_bb2_or163_i1732);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_9_i1129_stall_local;
wire local_bb2_reduction_9_i1129;

assign local_bb2_reduction_9_i1129 = (local_bb2_reduction_7_i1127 & local_bb2_reduction_8_i1128);

// This section implements an unregistered operation.
// 
wire local_bb2_or1237_i1168_stall_local;
wire [7:0] local_bb2_or1237_i1168;

assign local_bb2_or1237_i1168 = (local_bb2__30_i1162 | local_bb2__29_i1160);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i1170_stall_local;
wire [7:0] local_bb2__33_i1170;

assign local_bb2__33_i1170 = (local_bb2_cmp116_i1167 ? local_bb2__29_i1160 : local_bb2__31_i1164);

// This section implements an unregistered operation.
// 
wire local_bb2_or162_i1183_stall_local;
wire [31:0] local_bb2_or162_i1183;

assign local_bb2_or162_i1183 = (local_bb2_or1596_i1182 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_9_i117_stall_local;
wire local_bb2_reduction_9_i117;

assign local_bb2_reduction_9_i117 = (local_bb2_reduction_7_i115 & local_bb2_reduction_8_i116);

// This section implements an unregistered operation.
// 
wire local_bb2_or1237_i156_stall_local;
wire [7:0] local_bb2_or1237_i156;

assign local_bb2_or1237_i156 = (local_bb2__30_i150 | local_bb2__29_i148);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i158_stall_local;
wire [7:0] local_bb2__33_i158;

assign local_bb2__33_i158 = (local_bb2_cmp116_i155 ? local_bb2__29_i148 : local_bb2__31_i152);

// This section implements an unregistered operation.
// 
wire local_bb2_or162_i171_stall_local;
wire [31:0] local_bb2_or162_i171;

assign local_bb2_or162_i171 = (local_bb2_or1596_i170 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__26_i665_stall_local;
wire local_bb2__26_i665;

assign local_bb2__26_i665 = (local_bb2_reduction_9_i664 ? local_bb2_cmp38_i : local_bb2__24_i660);

// This section implements an unregistered operation.
// 
wire local_bb2_or124_i680_stall_local;
wire [31:0] local_bb2_or124_i680;

assign local_bb2_or124_i680[31:8] = 24'h0;
assign local_bb2_or124_i680[7:0] = local_bb2_or1247_i;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u121_stall_local;
wire [7:0] local_bb2_var__u121;

assign local_bb2_var__u121 = (local_bb2__33_i681 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__37_v_i684_stall_local;
wire [31:0] local_bb2__37_v_i684;

assign local_bb2__37_v_i684 = (local_bb2_Pivot20_i682 ? 32'h0 : local_bb2_or163_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or125_i1720_stall_local;
wire [31:0] local_bb2_or125_i1720;

assign local_bb2_or125_i1720 = (local_bb2_cmp117_i1716 ? 32'h0 : local_bb2_or124_i1718);

// This section implements an unregistered operation.
// 
wire local_bb2_conv136_i1722_stall_local;
wire [31:0] local_bb2_conv136_i1722;

assign local_bb2_conv136_i1722[31:8] = 24'h0;
assign local_bb2_conv136_i1722[7:0] = local_bb2_var__u120;

// This section implements an unregistered operation.
// 
wire local_bb2__39_v_i1734_stall_local;
wire [31:0] local_bb2__39_v_i1734;

assign local_bb2__39_v_i1734 = (local_bb2_SwitchLeaf_i1729 ? local_bb2_var__u104 : local_bb2__37_v_i1733);

// This section implements an unregistered operation.
// 
wire local_bb2__26_i1130_stall_local;
wire local_bb2__26_i1130;

assign local_bb2__26_i1130 = (local_bb2_reduction_9_i1129 ? local_bb2_cmp37_i1117 : local_bb2__24_i1125);

// This section implements an unregistered operation.
// 
wire local_bb2_or123_i1169_stall_local;
wire [31:0] local_bb2_or123_i1169;

assign local_bb2_or123_i1169[31:8] = 24'h0;
assign local_bb2_or123_i1169[7:0] = local_bb2_or1237_i1168;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u122_stall_local;
wire [7:0] local_bb2_var__u122;

assign local_bb2_var__u122 = (local_bb2__33_i1170 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__37_v_i1184_stall_local;
wire [31:0] local_bb2__37_v_i1184;

assign local_bb2__37_v_i1184 = (local_bb2_Pivot20_i1179 ? 32'h0 : local_bb2_or162_i1183);

// This section implements an unregistered operation.
// 
wire local_bb2__26_i118_stall_local;
wire local_bb2__26_i118;

assign local_bb2__26_i118 = (local_bb2_reduction_9_i117 ? local_bb2_cmp37_i105 : local_bb2__24_i113);

// This section implements an unregistered operation.
// 
wire local_bb2_or123_i157_stall_local;
wire [31:0] local_bb2_or123_i157;

assign local_bb2_or123_i157[31:8] = 24'h0;
assign local_bb2_or123_i157[7:0] = local_bb2_or1237_i156;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u123_stall_local;
wire [7:0] local_bb2_var__u123;

assign local_bb2_var__u123 = (local_bb2__33_i158 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__37_v_i172_stall_local;
wire [31:0] local_bb2__37_v_i172;

assign local_bb2__37_v_i172 = (local_bb2_Pivot20_i167 ? 32'h0 : local_bb2_or162_i171);

// This section implements an unregistered operation.
// 
wire local_bb2_or125_i_stall_local;
wire [31:0] local_bb2_or125_i;

assign local_bb2_or125_i = (local_bb2_cmp117_i ? 32'h0 : local_bb2_or124_i680);

// This section implements an unregistered operation.
// 
wire local_bb2_conv136_i_stall_local;
wire [31:0] local_bb2_conv136_i;

assign local_bb2_conv136_i[31:8] = 24'h0;
assign local_bb2_conv136_i[7:0] = local_bb2_var__u121;

// This section implements an unregistered operation.
// 
wire local_bb2__39_v_i685_stall_local;
wire [31:0] local_bb2__39_v_i685;

assign local_bb2__39_v_i685 = (local_bb2_SwitchLeaf_i683 ? local_bb2_var__u109 : local_bb2__37_v_i684);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i1735_stall_local;
wire [31:0] local_bb2_reduction_3_i1735;

assign local_bb2_reduction_3_i1735 = (local_bb2__32_i1714 | local_bb2_or125_i1720);

// This section implements an unregistered operation.
// 
wire local_bb2_or137_i1724_stall_local;
wire [31:0] local_bb2_or137_i1724;

assign local_bb2_or137_i1724 = (local_bb2_cmp132_not_i1723 ? local_bb2_conv136_i1722 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or124_i1171_stall_local;
wire [31:0] local_bb2_or124_i1171;

assign local_bb2_or124_i1171 = (local_bb2_cmp116_i1167 ? 32'h0 : local_bb2_or123_i1169);

// This section implements an unregistered operation.
// 
wire local_bb2_conv135_i1173_stall_local;
wire [31:0] local_bb2_conv135_i1173;

assign local_bb2_conv135_i1173[31:8] = 24'h0;
assign local_bb2_conv135_i1173[7:0] = local_bb2_var__u122;

// This section implements an unregistered operation.
// 
wire local_bb2__39_v_i1185_stall_local;
wire [31:0] local_bb2__39_v_i1185;

assign local_bb2__39_v_i1185 = (local_bb2_SwitchLeaf_i1180 ? local_bb2_var__u113 : local_bb2__37_v_i1184);

// This section implements an unregistered operation.
// 
wire local_bb2_or124_i159_stall_local;
wire [31:0] local_bb2_or124_i159;

assign local_bb2_or124_i159 = (local_bb2_cmp116_i155 ? 32'h0 : local_bb2_or123_i157);

// This section implements an unregistered operation.
// 
wire local_bb2_conv135_i161_stall_local;
wire [31:0] local_bb2_conv135_i161;

assign local_bb2_conv135_i161[31:8] = 24'h0;
assign local_bb2_conv135_i161[7:0] = local_bb2_var__u123;

// This section implements an unregistered operation.
// 
wire local_bb2__39_v_i173_stall_local;
wire [31:0] local_bb2__39_v_i173;

assign local_bb2__39_v_i173 = (local_bb2_SwitchLeaf_i168 ? local_bb2_var__u116 : local_bb2__37_v_i172);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i686_stall_local;
wire [31:0] local_bb2_reduction_3_i686;

assign local_bb2_reduction_3_i686 = (local_bb2__32_i679 | local_bb2_or125_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or137_i_stall_local;
wire [31:0] local_bb2_or137_i;

assign local_bb2_or137_i = (local_bb2_cmp132_not_i ? local_bb2_conv136_i : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i1737_stall_local;
wire [31:0] local_bb2_reduction_5_i1737;

assign local_bb2_reduction_5_i1737 = (local_bb2_shr151_i1727 | local_bb2_reduction_3_i1735);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_4_i1736_stall_local;
wire [31:0] local_bb2_reduction_4_i1736;

assign local_bb2_reduction_4_i1736 = (local_bb2_or137_i1724 | local_bb2__39_v_i1734);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i1186_stall_local;
wire [31:0] local_bb2_reduction_3_i1186;

assign local_bb2_reduction_3_i1186 = (local_bb2__32_i1165 | local_bb2_or124_i1171);

// This section implements an unregistered operation.
// 
wire local_bb2_or136_i1175_stall_local;
wire [31:0] local_bb2_or136_i1175;

assign local_bb2_or136_i1175 = (local_bb2_cmp131_not_i1174 ? local_bb2_conv135_i1173 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i174_stall_local;
wire [31:0] local_bb2_reduction_3_i174;

assign local_bb2_reduction_3_i174 = (local_bb2__32_i153 | local_bb2_or124_i159);

// This section implements an unregistered operation.
// 
wire local_bb2_or136_i163_stall_local;
wire [31:0] local_bb2_or136_i163;

assign local_bb2_or136_i163 = (local_bb2_cmp131_not_i162 ? local_bb2_conv135_i161 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i688_stall_local;
wire [31:0] local_bb2_reduction_5_i688;

assign local_bb2_reduction_5_i688 = (local_bb2_shr151_i | local_bb2_reduction_3_i686);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_4_i687_stall_local;
wire [31:0] local_bb2_reduction_4_i687;

assign local_bb2_reduction_4_i687 = (local_bb2_or137_i | local_bb2__39_v_i685);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i1738_stall_local;
wire [31:0] local_bb2_reduction_6_i1738;

assign local_bb2_reduction_6_i1738 = (local_bb2_reduction_4_i1736 | local_bb2_reduction_5_i1737);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i1188_stall_local;
wire [31:0] local_bb2_reduction_5_i1188;

assign local_bb2_reduction_5_i1188 = (local_bb2_shr150_i1178 | local_bb2_reduction_3_i1186);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_4_i1187_stall_local;
wire [31:0] local_bb2_reduction_4_i1187;

assign local_bb2_reduction_4_i1187 = (local_bb2_or136_i1175 | local_bb2__39_v_i1185);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i176_stall_local;
wire [31:0] local_bb2_reduction_5_i176;

assign local_bb2_reduction_5_i176 = (local_bb2_shr150_i166 | local_bb2_reduction_3_i174);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_4_i175_stall_local;
wire [31:0] local_bb2_reduction_4_i175;

assign local_bb2_reduction_4_i175 = (local_bb2_or136_i163 | local_bb2__39_v_i173);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i689_stall_local;
wire [31:0] local_bb2_reduction_6_i689;

assign local_bb2_reduction_6_i689 = (local_bb2_reduction_4_i687 | local_bb2_reduction_5_i688);

// This section implements an unregistered operation.
// 
wire local_bb2_xor189_i1740_stall_local;
wire [31:0] local_bb2_xor189_i1740;

assign local_bb2_xor189_i1740 = (local_bb2_reduction_6_i1738 ^ local_bb2_xor36_lobit_i1739);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i1189_stall_local;
wire [31:0] local_bb2_reduction_6_i1189;

assign local_bb2_reduction_6_i1189 = (local_bb2_reduction_4_i1187 | local_bb2_reduction_5_i1188);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i177_stall_local;
wire [31:0] local_bb2_reduction_6_i177;

assign local_bb2_reduction_6_i177 = (local_bb2_reduction_4_i175 | local_bb2_reduction_5_i176);

// This section implements an unregistered operation.
// 
wire local_bb2_xor189_i_stall_local;
wire [31:0] local_bb2_xor189_i;

assign local_bb2_xor189_i = (local_bb2_reduction_6_i689 ^ local_bb2_xor36_lobit_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp38_i1666_valid_out_1;
wire local_bb2_cmp38_i1666_stall_in_1;
 reg local_bb2_cmp38_i1666_consumed_1_NO_SHIFT_REG;
wire local_bb2__26_i1679_valid_out;
wire local_bb2__26_i1679_stall_in;
 reg local_bb2__26_i1679_consumed_0_NO_SHIFT_REG;
wire local_bb2_add193_i1743_valid_out;
wire local_bb2_add193_i1743_stall_in;
 reg local_bb2_add193_i1743_consumed_0_NO_SHIFT_REG;
wire local_bb2_and17_i1655_valid_out_2;
wire local_bb2_and17_i1655_stall_in_2;
 reg local_bb2_and17_i1655_consumed_2_NO_SHIFT_REG;
wire local_bb2_var__u102_valid_out;
wire local_bb2_var__u102_stall_in;
 reg local_bb2_var__u102_consumed_0_NO_SHIFT_REG;
wire local_bb2_add193_i1743_inputs_ready;
wire local_bb2_add193_i1743_stall_local;
wire [31:0] local_bb2_add193_i1743;

assign local_bb2_add193_i1743_inputs_ready = (rnode_172to173_bb2__22_i1652_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i1663_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_lnot23_i1661_0_valid_out_NO_SHIFT_REG & rnode_172to173_bb2__22_i1652_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2__23_i1653_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2__23_i1653_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i1663_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2_shr16_i1654_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i1663_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1689_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1689_0_valid_out_4_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1689_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1689_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1689_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_add193_i1743 = (local_bb2_add_i1742 + local_bb2_xor189_i1740);
assign local_bb2_cmp38_i1666_valid_out_1 = 1'b1;
assign local_bb2__26_i1679_valid_out = 1'b1;
assign local_bb2_add193_i1743_valid_out = 1'b1;
assign local_bb2_and17_i1655_valid_out_2 = 1'b1;
assign local_bb2_var__u102_valid_out = 1'b1;
assign rnode_172to173_bb2__22_i1652_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i1663_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_lnot23_i1661_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i1652_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i1653_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i1653_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i1663_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_shr16_i1654_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i1663_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1689_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1689_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1689_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1689_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1689_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp38_i1666_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__26_i1679_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add193_i1743_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and17_i1655_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u102_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp38_i1666_consumed_1_NO_SHIFT_REG <= (local_bb2_add193_i1743_inputs_ready & (local_bb2_cmp38_i1666_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp38_i1666_stall_in_1)) & local_bb2_add193_i1743_stall_local);
		local_bb2__26_i1679_consumed_0_NO_SHIFT_REG <= (local_bb2_add193_i1743_inputs_ready & (local_bb2__26_i1679_consumed_0_NO_SHIFT_REG | ~(local_bb2__26_i1679_stall_in)) & local_bb2_add193_i1743_stall_local);
		local_bb2_add193_i1743_consumed_0_NO_SHIFT_REG <= (local_bb2_add193_i1743_inputs_ready & (local_bb2_add193_i1743_consumed_0_NO_SHIFT_REG | ~(local_bb2_add193_i1743_stall_in)) & local_bb2_add193_i1743_stall_local);
		local_bb2_and17_i1655_consumed_2_NO_SHIFT_REG <= (local_bb2_add193_i1743_inputs_ready & (local_bb2_and17_i1655_consumed_2_NO_SHIFT_REG | ~(local_bb2_and17_i1655_stall_in_2)) & local_bb2_add193_i1743_stall_local);
		local_bb2_var__u102_consumed_0_NO_SHIFT_REG <= (local_bb2_add193_i1743_inputs_ready & (local_bb2_var__u102_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u102_stall_in)) & local_bb2_add193_i1743_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_xor188_i1191_stall_local;
wire [31:0] local_bb2_xor188_i1191;

assign local_bb2_xor188_i1191 = (local_bb2_reduction_6_i1189 ^ local_bb2_xor_lobit_i1190);

// This section implements an unregistered operation.
// 
wire local_bb2_xor188_i179_stall_local;
wire [31:0] local_bb2_xor188_i179;

assign local_bb2_xor188_i179 = (local_bb2_reduction_6_i177 ^ local_bb2_xor_lobit_i178);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp38_i_valid_out_1;
wire local_bb2_cmp38_i_stall_in_1;
 reg local_bb2_cmp38_i_consumed_1_NO_SHIFT_REG;
wire local_bb2__26_i665_valid_out;
wire local_bb2__26_i665_stall_in;
 reg local_bb2__26_i665_consumed_0_NO_SHIFT_REG;
wire local_bb2_add193_i_valid_out;
wire local_bb2_add193_i_stall_in;
 reg local_bb2_add193_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_and17_i643_valid_out_2;
wire local_bb2_and17_i643_stall_in_2;
 reg local_bb2_and17_i643_consumed_2_NO_SHIFT_REG;
wire local_bb2_var__u107_valid_out;
wire local_bb2_var__u107_stall_in;
 reg local_bb2_var__u107_consumed_0_NO_SHIFT_REG;
wire local_bb2_add193_i_inputs_ready;
wire local_bb2_add193_i_stall_local;
wire [31:0] local_bb2_add193_i;

assign local_bb2_add193_i_inputs_ready = (rnode_172to173_bb2__22_i640_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i651_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_lnot23_i649_0_valid_out_NO_SHIFT_REG & rnode_172to173_bb2__22_i640_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2__23_i641_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2__23_i641_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i651_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2_shr16_i642_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i651_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i671_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i671_0_valid_out_4_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i671_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i671_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i671_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_add193_i = (local_bb2_add_i690 + local_bb2_xor189_i);
assign local_bb2_cmp38_i_valid_out_1 = 1'b1;
assign local_bb2__26_i665_valid_out = 1'b1;
assign local_bb2_add193_i_valid_out = 1'b1;
assign local_bb2_and17_i643_valid_out_2 = 1'b1;
assign local_bb2_var__u107_valid_out = 1'b1;
assign rnode_172to173_bb2__22_i640_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i651_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_lnot23_i649_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i640_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i641_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i641_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i651_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_shr16_i642_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i651_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i671_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i671_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i671_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i671_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i671_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp38_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__26_i665_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add193_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and17_i643_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u107_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp38_i_consumed_1_NO_SHIFT_REG <= (local_bb2_add193_i_inputs_ready & (local_bb2_cmp38_i_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp38_i_stall_in_1)) & local_bb2_add193_i_stall_local);
		local_bb2__26_i665_consumed_0_NO_SHIFT_REG <= (local_bb2_add193_i_inputs_ready & (local_bb2__26_i665_consumed_0_NO_SHIFT_REG | ~(local_bb2__26_i665_stall_in)) & local_bb2_add193_i_stall_local);
		local_bb2_add193_i_consumed_0_NO_SHIFT_REG <= (local_bb2_add193_i_inputs_ready & (local_bb2_add193_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_add193_i_stall_in)) & local_bb2_add193_i_stall_local);
		local_bb2_and17_i643_consumed_2_NO_SHIFT_REG <= (local_bb2_add193_i_inputs_ready & (local_bb2_and17_i643_consumed_2_NO_SHIFT_REG | ~(local_bb2_and17_i643_stall_in_2)) & local_bb2_add193_i_stall_local);
		local_bb2_var__u107_consumed_0_NO_SHIFT_REG <= (local_bb2_add193_i_inputs_ready & (local_bb2_var__u107_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u107_stall_in)) & local_bb2_add193_i_stall_local);
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_cmp38_i1666_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i1666_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_cmp38_i1666_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_cmp38_i1666_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_cmp38_i1666_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_cmp38_i1666_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_cmp38_i1666_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_cmp38_i1666),
	.data_out(rnode_173to175_bb2_cmp38_i1666_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_cmp38_i1666_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_cmp38_i1666_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_173to175_bb2_cmp38_i1666_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_cmp38_i1666_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_cmp38_i1666_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp38_i1666_stall_in_1 = 1'b0;
assign rnode_173to175_bb2_cmp38_i1666_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp38_i1666_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp38_i1666_0_NO_SHIFT_REG = rnode_173to175_bb2_cmp38_i1666_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_cmp38_i1666_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp38_i1666_1_NO_SHIFT_REG = rnode_173to175_bb2_cmp38_i1666_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_cmp38_i1666_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp38_i1666_2_NO_SHIFT_REG = rnode_173to175_bb2_cmp38_i1666_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2__26_i1679_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1679_0_stall_in_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1679_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1679_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1679_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1679_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1679_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1679_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2__26_i1679_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2__26_i1679_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2__26_i1679_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2__26_i1679_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2__26_i1679_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2__26_i1679),
	.data_out(rnode_173to174_bb2__26_i1679_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2__26_i1679_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2__26_i1679_0_reg_174_fifo.DATA_WIDTH = 1;
defparam rnode_173to174_bb2__26_i1679_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2__26_i1679_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2__26_i1679_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__26_i1679_stall_in = 1'b0;
assign rnode_173to174_bb2__26_i1679_0_NO_SHIFT_REG = rnode_173to174_bb2__26_i1679_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2__26_i1679_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2__26_i1679_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_add193_i1743_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i1743_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i1743_1_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i1743_2_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i1743_3_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i1743_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_valid_out_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_stall_in_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i1743_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_add193_i1743_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_add193_i1743_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_add193_i1743_0_stall_in_0_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_add193_i1743_0_valid_out_0_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_add193_i1743_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_add193_i1743),
	.data_out(rnode_173to174_bb2_add193_i1743_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_add193_i1743_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_add193_i1743_0_reg_174_fifo.DATA_WIDTH = 32;
defparam rnode_173to174_bb2_add193_i1743_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_add193_i1743_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_add193_i1743_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add193_i1743_stall_in = 1'b0;
assign rnode_173to174_bb2_add193_i1743_0_stall_in_0_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_add193_i1743_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add193_i1743_0_NO_SHIFT_REG = rnode_173to174_bb2_add193_i1743_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add193_i1743_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add193_i1743_1_NO_SHIFT_REG = rnode_173to174_bb2_add193_i1743_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add193_i1743_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add193_i1743_2_NO_SHIFT_REG = rnode_173to174_bb2_add193_i1743_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add193_i1743_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add193_i1743_3_NO_SHIFT_REG = rnode_173to174_bb2_add193_i1743_0_reg_174_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_and17_i1655_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1655_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_and17_i1655_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1655_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_and17_i1655_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1655_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1655_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1655_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_and17_i1655_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_and17_i1655_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_and17_i1655_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_and17_i1655_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_and17_i1655_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and17_i1655),
	.data_out(rnode_173to175_bb2_and17_i1655_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_and17_i1655_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_and17_i1655_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_173to175_bb2_and17_i1655_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_and17_i1655_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_and17_i1655_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and17_i1655_stall_in_2 = 1'b0;
assign rnode_173to175_bb2_and17_i1655_0_NO_SHIFT_REG = rnode_173to175_bb2_and17_i1655_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_and17_i1655_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_and17_i1655_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_var__u102_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u102_0_stall_in_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u102_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u102_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u102_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u102_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u102_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u102_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_var__u102_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_var__u102_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_var__u102_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_var__u102_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_var__u102_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_var__u102),
	.data_out(rnode_173to174_bb2_var__u102_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_var__u102_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_var__u102_0_reg_174_fifo.DATA_WIDTH = 1;
defparam rnode_173to174_bb2_var__u102_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_var__u102_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_var__u102_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u102_stall_in = 1'b0;
assign rnode_173to174_bb2_var__u102_0_NO_SHIFT_REG = rnode_173to174_bb2_var__u102_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_var__u102_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_var__u102_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i1117_valid_out_1;
wire local_bb2_cmp37_i1117_stall_in_1;
 reg local_bb2_cmp37_i1117_consumed_1_NO_SHIFT_REG;
wire local_bb2__26_i1130_valid_out;
wire local_bb2__26_i1130_stall_in;
 reg local_bb2__26_i1130_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i1194_valid_out;
wire local_bb2_add192_i1194_stall_in;
 reg local_bb2_add192_i1194_consumed_0_NO_SHIFT_REG;
wire local_bb2_and17_i1106_valid_out_2;
wire local_bb2_and17_i1106_stall_in_2;
 reg local_bb2_and17_i1106_consumed_2_NO_SHIFT_REG;
wire local_bb2_var__u111_valid_out;
wire local_bb2_var__u111_stall_in;
 reg local_bb2_var__u111_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i1194_inputs_ready;
wire local_bb2_add192_i1194_stall_local;
wire [31:0] local_bb2_add192_i1194;

assign local_bb2_add192_i1194_inputs_ready = (rnode_172to173_bb2__22_i1103_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i1114_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_lnot23_i1112_0_valid_out_NO_SHIFT_REG & rnode_172to173_bb2__22_i1103_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2__23_i1104_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2__23_i1104_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i1114_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2_shr16_i1105_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i1114_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1140_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1140_0_valid_out_4_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1140_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1140_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i1140_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_add192_i1194 = (local_bb2_add_i1193 + local_bb2_xor188_i1191);
assign local_bb2_cmp37_i1117_valid_out_1 = 1'b1;
assign local_bb2__26_i1130_valid_out = 1'b1;
assign local_bb2_add192_i1194_valid_out = 1'b1;
assign local_bb2_and17_i1106_valid_out_2 = 1'b1;
assign local_bb2_var__u111_valid_out = 1'b1;
assign rnode_172to173_bb2__22_i1103_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i1114_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_lnot23_i1112_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i1103_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i1104_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i1104_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i1114_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_shr16_i1105_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i1114_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1140_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1140_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1140_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1140_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i1140_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp37_i1117_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__26_i1130_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add192_i1194_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and17_i1106_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u111_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp37_i1117_consumed_1_NO_SHIFT_REG <= (local_bb2_add192_i1194_inputs_ready & (local_bb2_cmp37_i1117_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp37_i1117_stall_in_1)) & local_bb2_add192_i1194_stall_local);
		local_bb2__26_i1130_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1194_inputs_ready & (local_bb2__26_i1130_consumed_0_NO_SHIFT_REG | ~(local_bb2__26_i1130_stall_in)) & local_bb2_add192_i1194_stall_local);
		local_bb2_add192_i1194_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1194_inputs_ready & (local_bb2_add192_i1194_consumed_0_NO_SHIFT_REG | ~(local_bb2_add192_i1194_stall_in)) & local_bb2_add192_i1194_stall_local);
		local_bb2_and17_i1106_consumed_2_NO_SHIFT_REG <= (local_bb2_add192_i1194_inputs_ready & (local_bb2_and17_i1106_consumed_2_NO_SHIFT_REG | ~(local_bb2_and17_i1106_stall_in_2)) & local_bb2_add192_i1194_stall_local);
		local_bb2_var__u111_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1194_inputs_ready & (local_bb2_var__u111_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u111_stall_in)) & local_bb2_add192_i1194_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i105_valid_out_1;
wire local_bb2_cmp37_i105_stall_in_1;
 reg local_bb2_cmp37_i105_consumed_1_NO_SHIFT_REG;
wire local_bb2__26_i118_valid_out;
wire local_bb2__26_i118_stall_in;
 reg local_bb2__26_i118_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i182_valid_out;
wire local_bb2_add192_i182_stall_in;
 reg local_bb2_add192_i182_consumed_0_NO_SHIFT_REG;
wire local_bb2_and17_i94_valid_out_2;
wire local_bb2_and17_i94_stall_in_2;
 reg local_bb2_and17_i94_consumed_2_NO_SHIFT_REG;
wire local_bb2_var__u114_valid_out;
wire local_bb2_var__u114_stall_in;
 reg local_bb2_var__u114_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i182_inputs_ready;
wire local_bb2_add192_i182_stall_local;
wire [31:0] local_bb2_add192_i182;

assign local_bb2_add192_i182_inputs_ready = (rnode_172to173_bb2__22_i91_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i102_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_lnot23_i100_0_valid_out_NO_SHIFT_REG & rnode_172to173_bb2__22_i91_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2__23_i92_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2__23_i92_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i102_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2_shr16_i93_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_cmp27_i102_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i128_0_valid_out_0_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i128_0_valid_out_4_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i128_0_valid_out_1_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i128_0_valid_out_2_NO_SHIFT_REG & rnode_172to173_bb2_align_0_i128_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_add192_i182 = (local_bb2_add_i181 + local_bb2_xor188_i179);
assign local_bb2_cmp37_i105_valid_out_1 = 1'b1;
assign local_bb2__26_i118_valid_out = 1'b1;
assign local_bb2_add192_i182_valid_out = 1'b1;
assign local_bb2_and17_i94_valid_out_2 = 1'b1;
assign local_bb2_var__u114_valid_out = 1'b1;
assign rnode_172to173_bb2__22_i91_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i102_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_lnot23_i100_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__22_i91_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i92_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2__23_i92_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i102_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_shr16_i93_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_cmp27_i102_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i128_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i128_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i128_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i128_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_172to173_bb2_align_0_i128_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp37_i105_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__26_i118_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add192_i182_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and17_i94_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u114_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp37_i105_consumed_1_NO_SHIFT_REG <= (local_bb2_add192_i182_inputs_ready & (local_bb2_cmp37_i105_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp37_i105_stall_in_1)) & local_bb2_add192_i182_stall_local);
		local_bb2__26_i118_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i182_inputs_ready & (local_bb2__26_i118_consumed_0_NO_SHIFT_REG | ~(local_bb2__26_i118_stall_in)) & local_bb2_add192_i182_stall_local);
		local_bb2_add192_i182_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i182_inputs_ready & (local_bb2_add192_i182_consumed_0_NO_SHIFT_REG | ~(local_bb2_add192_i182_stall_in)) & local_bb2_add192_i182_stall_local);
		local_bb2_and17_i94_consumed_2_NO_SHIFT_REG <= (local_bb2_add192_i182_inputs_ready & (local_bb2_and17_i94_consumed_2_NO_SHIFT_REG | ~(local_bb2_and17_i94_stall_in_2)) & local_bb2_add192_i182_stall_local);
		local_bb2_var__u114_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i182_inputs_ready & (local_bb2_var__u114_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u114_stall_in)) & local_bb2_add192_i182_stall_local);
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_cmp38_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp38_i_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_cmp38_i_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_cmp38_i_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_cmp38_i_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_cmp38_i_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_cmp38_i_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_cmp38_i),
	.data_out(rnode_173to175_bb2_cmp38_i_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_cmp38_i_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_cmp38_i_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_173to175_bb2_cmp38_i_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_cmp38_i_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_cmp38_i_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp38_i_stall_in_1 = 1'b0;
assign rnode_173to175_bb2_cmp38_i_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp38_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp38_i_0_NO_SHIFT_REG = rnode_173to175_bb2_cmp38_i_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_cmp38_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp38_i_1_NO_SHIFT_REG = rnode_173to175_bb2_cmp38_i_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_cmp38_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp38_i_2_NO_SHIFT_REG = rnode_173to175_bb2_cmp38_i_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2__26_i665_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i665_0_stall_in_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i665_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i665_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i665_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i665_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i665_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i665_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2__26_i665_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2__26_i665_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2__26_i665_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2__26_i665_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2__26_i665_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2__26_i665),
	.data_out(rnode_173to174_bb2__26_i665_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2__26_i665_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2__26_i665_0_reg_174_fifo.DATA_WIDTH = 1;
defparam rnode_173to174_bb2__26_i665_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2__26_i665_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2__26_i665_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__26_i665_stall_in = 1'b0;
assign rnode_173to174_bb2__26_i665_0_NO_SHIFT_REG = rnode_173to174_bb2__26_i665_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2__26_i665_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2__26_i665_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_add193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i_1_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i_2_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i_3_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add193_i_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_valid_out_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_stall_in_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add193_i_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_add193_i_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_add193_i_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_add193_i_0_stall_in_0_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_add193_i_0_valid_out_0_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_add193_i_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_add193_i),
	.data_out(rnode_173to174_bb2_add193_i_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_add193_i_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_add193_i_0_reg_174_fifo.DATA_WIDTH = 32;
defparam rnode_173to174_bb2_add193_i_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_add193_i_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_add193_i_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add193_i_stall_in = 1'b0;
assign rnode_173to174_bb2_add193_i_0_stall_in_0_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_add193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add193_i_0_NO_SHIFT_REG = rnode_173to174_bb2_add193_i_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add193_i_1_NO_SHIFT_REG = rnode_173to174_bb2_add193_i_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add193_i_2_NO_SHIFT_REG = rnode_173to174_bb2_add193_i_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add193_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add193_i_3_NO_SHIFT_REG = rnode_173to174_bb2_add193_i_0_reg_174_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_and17_i643_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i643_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_and17_i643_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i643_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_and17_i643_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i643_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i643_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i643_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_and17_i643_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_and17_i643_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_and17_i643_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_and17_i643_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_and17_i643_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and17_i643),
	.data_out(rnode_173to175_bb2_and17_i643_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_and17_i643_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_and17_i643_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_173to175_bb2_and17_i643_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_and17_i643_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_and17_i643_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and17_i643_stall_in_2 = 1'b0;
assign rnode_173to175_bb2_and17_i643_0_NO_SHIFT_REG = rnode_173to175_bb2_and17_i643_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_and17_i643_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_and17_i643_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_var__u107_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u107_0_stall_in_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u107_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u107_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u107_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u107_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u107_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u107_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_var__u107_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_var__u107_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_var__u107_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_var__u107_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_var__u107_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_var__u107),
	.data_out(rnode_173to174_bb2_var__u107_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_var__u107_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_var__u107_0_reg_174_fifo.DATA_WIDTH = 1;
defparam rnode_173to174_bb2_var__u107_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_var__u107_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_var__u107_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u107_stall_in = 1'b0;
assign rnode_173to174_bb2_var__u107_0_NO_SHIFT_REG = rnode_173to174_bb2_var__u107_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_var__u107_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_var__u107_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_not_cmp38_i1772_stall_local;
wire local_bb2_not_cmp38_i1772;

assign local_bb2_not_cmp38_i1772 = (rnode_173to175_bb2_cmp38_i1666_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2__26_i1679_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1679_0_stall_in_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1679_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1679_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1679_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1679_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1679_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1679_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2__26_i1679_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2__26_i1679_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2__26_i1679_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2__26_i1679_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2__26_i1679_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2__26_i1679_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2__26_i1679_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2__26_i1679_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2__26_i1679_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_174to175_bb2__26_i1679_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2__26_i1679_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2__26_i1679_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2__26_i1679_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__26_i1679_0_NO_SHIFT_REG = rnode_174to175_bb2__26_i1679_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__26_i1679_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__26_i1679_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and194_i1744_valid_out;
wire local_bb2_and194_i1744_stall_in;
wire local_bb2_and194_i1744_inputs_ready;
wire local_bb2_and194_i1744_stall_local;
wire [31:0] local_bb2_and194_i1744;

assign local_bb2_and194_i1744_inputs_ready = rnode_173to174_bb2_add193_i1743_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_and194_i1744 = (rnode_173to174_bb2_add193_i1743_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb2_and194_i1744_valid_out = 1'b1;
assign rnode_173to174_bb2_add193_i1743_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and196_i1745_valid_out;
wire local_bb2_and196_i1745_stall_in;
wire local_bb2_and196_i1745_inputs_ready;
wire local_bb2_and196_i1745_stall_local;
wire [31:0] local_bb2_and196_i1745;

assign local_bb2_and196_i1745_inputs_ready = rnode_173to174_bb2_add193_i1743_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and196_i1745 = (rnode_173to174_bb2_add193_i1743_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb2_and196_i1745_valid_out = 1'b1;
assign rnode_173to174_bb2_add193_i1743_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and199_i1746_valid_out;
wire local_bb2_and199_i1746_stall_in;
wire local_bb2_and199_i1746_inputs_ready;
wire local_bb2_and199_i1746_stall_local;
wire [31:0] local_bb2_and199_i1746;

assign local_bb2_and199_i1746_inputs_ready = rnode_173to174_bb2_add193_i1743_0_valid_out_2_NO_SHIFT_REG;
assign local_bb2_and199_i1746 = (rnode_173to174_bb2_add193_i1743_2_NO_SHIFT_REG & 32'h1);
assign local_bb2_and199_i1746_valid_out = 1'b1;
assign rnode_173to174_bb2_add193_i1743_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and202_i1747_stall_local;
wire [31:0] local_bb2_and202_i1747;

assign local_bb2_and202_i1747 = (rnode_173to174_bb2_add193_i1743_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_var__u102_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u102_0_stall_in_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u102_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u102_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u102_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u102_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u102_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u102_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_var__u102_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_var__u102_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_var__u102_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_var__u102_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_var__u102_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2_var__u102_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2_var__u102_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_var__u102_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_var__u102_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_174to175_bb2_var__u102_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_var__u102_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_var__u102_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_var__u102_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_var__u102_0_NO_SHIFT_REG = rnode_174to175_bb2_var__u102_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_var__u102_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_var__u102_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_cmp37_i1117_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i1117_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_cmp37_i1117_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_cmp37_i1117_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_cmp37_i1117_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_cmp37_i1117_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_cmp37_i1117_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_cmp37_i1117),
	.data_out(rnode_173to175_bb2_cmp37_i1117_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_cmp37_i1117_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_cmp37_i1117_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_173to175_bb2_cmp37_i1117_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_cmp37_i1117_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_cmp37_i1117_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp37_i1117_stall_in_1 = 1'b0;
assign rnode_173to175_bb2_cmp37_i1117_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp37_i1117_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp37_i1117_0_NO_SHIFT_REG = rnode_173to175_bb2_cmp37_i1117_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_cmp37_i1117_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp37_i1117_1_NO_SHIFT_REG = rnode_173to175_bb2_cmp37_i1117_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_cmp37_i1117_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp37_i1117_2_NO_SHIFT_REG = rnode_173to175_bb2_cmp37_i1117_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2__26_i1130_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1130_0_stall_in_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1130_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1130_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1130_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1130_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1130_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i1130_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2__26_i1130_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2__26_i1130_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2__26_i1130_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2__26_i1130_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2__26_i1130_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2__26_i1130),
	.data_out(rnode_173to174_bb2__26_i1130_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2__26_i1130_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2__26_i1130_0_reg_174_fifo.DATA_WIDTH = 1;
defparam rnode_173to174_bb2__26_i1130_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2__26_i1130_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2__26_i1130_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__26_i1130_stall_in = 1'b0;
assign rnode_173to174_bb2__26_i1130_0_NO_SHIFT_REG = rnode_173to174_bb2__26_i1130_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2__26_i1130_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2__26_i1130_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_add192_i1194_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i1194_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i1194_1_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i1194_2_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i1194_3_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i1194_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_valid_out_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_stall_in_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i1194_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_add192_i1194_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_add192_i1194_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_add192_i1194_0_stall_in_0_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_add192_i1194_0_valid_out_0_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_add192_i1194_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_add192_i1194),
	.data_out(rnode_173to174_bb2_add192_i1194_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_add192_i1194_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_add192_i1194_0_reg_174_fifo.DATA_WIDTH = 32;
defparam rnode_173to174_bb2_add192_i1194_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_add192_i1194_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_add192_i1194_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add192_i1194_stall_in = 1'b0;
assign rnode_173to174_bb2_add192_i1194_0_stall_in_0_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_add192_i1194_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add192_i1194_0_NO_SHIFT_REG = rnode_173to174_bb2_add192_i1194_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add192_i1194_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add192_i1194_1_NO_SHIFT_REG = rnode_173to174_bb2_add192_i1194_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add192_i1194_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add192_i1194_2_NO_SHIFT_REG = rnode_173to174_bb2_add192_i1194_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add192_i1194_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add192_i1194_3_NO_SHIFT_REG = rnode_173to174_bb2_add192_i1194_0_reg_174_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_and17_i1106_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1106_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_and17_i1106_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1106_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_and17_i1106_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1106_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1106_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i1106_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_and17_i1106_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_and17_i1106_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_and17_i1106_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_and17_i1106_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_and17_i1106_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and17_i1106),
	.data_out(rnode_173to175_bb2_and17_i1106_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_and17_i1106_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_and17_i1106_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_173to175_bb2_and17_i1106_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_and17_i1106_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_and17_i1106_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and17_i1106_stall_in_2 = 1'b0;
assign rnode_173to175_bb2_and17_i1106_0_NO_SHIFT_REG = rnode_173to175_bb2_and17_i1106_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_and17_i1106_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_and17_i1106_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_var__u111_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u111_0_stall_in_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u111_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u111_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u111_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u111_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u111_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u111_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_var__u111_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_var__u111_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_var__u111_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_var__u111_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_var__u111_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_var__u111),
	.data_out(rnode_173to174_bb2_var__u111_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_var__u111_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_var__u111_0_reg_174_fifo.DATA_WIDTH = 1;
defparam rnode_173to174_bb2_var__u111_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_var__u111_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_var__u111_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u111_stall_in = 1'b0;
assign rnode_173to174_bb2_var__u111_0_NO_SHIFT_REG = rnode_173to174_bb2_var__u111_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_var__u111_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_var__u111_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_cmp37_i105_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_1_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_2_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_cmp37_i105_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_cmp37_i105_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_cmp37_i105_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_cmp37_i105_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_cmp37_i105_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_cmp37_i105_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_cmp37_i105),
	.data_out(rnode_173to175_bb2_cmp37_i105_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_cmp37_i105_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_cmp37_i105_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_173to175_bb2_cmp37_i105_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_cmp37_i105_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_cmp37_i105_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp37_i105_stall_in_1 = 1'b0;
assign rnode_173to175_bb2_cmp37_i105_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp37_i105_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp37_i105_0_NO_SHIFT_REG = rnode_173to175_bb2_cmp37_i105_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_cmp37_i105_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp37_i105_1_NO_SHIFT_REG = rnode_173to175_bb2_cmp37_i105_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_cmp37_i105_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_173to175_bb2_cmp37_i105_2_NO_SHIFT_REG = rnode_173to175_bb2_cmp37_i105_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2__26_i118_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i118_0_stall_in_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i118_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i118_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i118_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i118_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i118_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2__26_i118_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2__26_i118_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2__26_i118_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2__26_i118_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2__26_i118_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2__26_i118_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2__26_i118),
	.data_out(rnode_173to174_bb2__26_i118_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2__26_i118_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2__26_i118_0_reg_174_fifo.DATA_WIDTH = 1;
defparam rnode_173to174_bb2__26_i118_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2__26_i118_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2__26_i118_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__26_i118_stall_in = 1'b0;
assign rnode_173to174_bb2__26_i118_0_NO_SHIFT_REG = rnode_173to174_bb2__26_i118_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2__26_i118_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2__26_i118_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_add192_i182_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i182_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i182_1_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i182_2_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i182_3_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to174_bb2_add192_i182_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_valid_out_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_stall_in_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_add192_i182_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_add192_i182_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_add192_i182_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_add192_i182_0_stall_in_0_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_add192_i182_0_valid_out_0_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_add192_i182_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_add192_i182),
	.data_out(rnode_173to174_bb2_add192_i182_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_add192_i182_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_add192_i182_0_reg_174_fifo.DATA_WIDTH = 32;
defparam rnode_173to174_bb2_add192_i182_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_add192_i182_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_add192_i182_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add192_i182_stall_in = 1'b0;
assign rnode_173to174_bb2_add192_i182_0_stall_in_0_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_add192_i182_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add192_i182_0_NO_SHIFT_REG = rnode_173to174_bb2_add192_i182_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add192_i182_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add192_i182_1_NO_SHIFT_REG = rnode_173to174_bb2_add192_i182_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add192_i182_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add192_i182_2_NO_SHIFT_REG = rnode_173to174_bb2_add192_i182_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_add192_i182_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_add192_i182_3_NO_SHIFT_REG = rnode_173to174_bb2_add192_i182_0_reg_174_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_173to175_bb2_and17_i94_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i94_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_and17_i94_0_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i94_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_173to175_bb2_and17_i94_0_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i94_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i94_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_173to175_bb2_and17_i94_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_173to175_bb2_and17_i94_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to175_bb2_and17_i94_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to175_bb2_and17_i94_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_173to175_bb2_and17_i94_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_173to175_bb2_and17_i94_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and17_i94),
	.data_out(rnode_173to175_bb2_and17_i94_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_173to175_bb2_and17_i94_0_reg_175_fifo.DEPTH = 2;
defparam rnode_173to175_bb2_and17_i94_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_173to175_bb2_and17_i94_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to175_bb2_and17_i94_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_173to175_bb2_and17_i94_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and17_i94_stall_in_2 = 1'b0;
assign rnode_173to175_bb2_and17_i94_0_NO_SHIFT_REG = rnode_173to175_bb2_and17_i94_0_reg_175_NO_SHIFT_REG;
assign rnode_173to175_bb2_and17_i94_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_and17_i94_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_173to174_bb2_var__u114_0_valid_out_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u114_0_stall_in_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u114_0_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u114_0_reg_174_inputs_ready_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u114_0_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u114_0_valid_out_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u114_0_stall_in_reg_174_NO_SHIFT_REG;
 logic rnode_173to174_bb2_var__u114_0_stall_out_reg_174_NO_SHIFT_REG;

acl_data_fifo rnode_173to174_bb2_var__u114_0_reg_174_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_173to174_bb2_var__u114_0_reg_174_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_173to174_bb2_var__u114_0_stall_in_reg_174_NO_SHIFT_REG),
	.valid_out(rnode_173to174_bb2_var__u114_0_valid_out_reg_174_NO_SHIFT_REG),
	.stall_out(rnode_173to174_bb2_var__u114_0_stall_out_reg_174_NO_SHIFT_REG),
	.data_in(local_bb2_var__u114),
	.data_out(rnode_173to174_bb2_var__u114_0_reg_174_NO_SHIFT_REG)
);

defparam rnode_173to174_bb2_var__u114_0_reg_174_fifo.DEPTH = 1;
defparam rnode_173to174_bb2_var__u114_0_reg_174_fifo.DATA_WIDTH = 1;
defparam rnode_173to174_bb2_var__u114_0_reg_174_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_173to174_bb2_var__u114_0_reg_174_fifo.IMPL = "shift_reg";

assign rnode_173to174_bb2_var__u114_0_reg_174_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u114_stall_in = 1'b0;
assign rnode_173to174_bb2_var__u114_0_NO_SHIFT_REG = rnode_173to174_bb2_var__u114_0_reg_174_NO_SHIFT_REG;
assign rnode_173to174_bb2_var__u114_0_stall_in_reg_174_NO_SHIFT_REG = 1'b0;
assign rnode_173to174_bb2_var__u114_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_not_cmp38_i_stall_local;
wire local_bb2_not_cmp38_i;

assign local_bb2_not_cmp38_i = (rnode_173to175_bb2_cmp38_i_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2__26_i665_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i665_0_stall_in_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i665_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i665_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i665_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i665_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i665_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i665_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2__26_i665_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2__26_i665_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2__26_i665_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2__26_i665_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2__26_i665_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2__26_i665_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2__26_i665_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2__26_i665_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2__26_i665_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_174to175_bb2__26_i665_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2__26_i665_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2__26_i665_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2__26_i665_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__26_i665_0_NO_SHIFT_REG = rnode_174to175_bb2__26_i665_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__26_i665_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__26_i665_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and194_i_valid_out;
wire local_bb2_and194_i_stall_in;
wire local_bb2_and194_i_inputs_ready;
wire local_bb2_and194_i_stall_local;
wire [31:0] local_bb2_and194_i;

assign local_bb2_and194_i_inputs_ready = rnode_173to174_bb2_add193_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_and194_i = (rnode_173to174_bb2_add193_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb2_and194_i_valid_out = 1'b1;
assign rnode_173to174_bb2_add193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and196_i_valid_out;
wire local_bb2_and196_i_stall_in;
wire local_bb2_and196_i_inputs_ready;
wire local_bb2_and196_i_stall_local;
wire [31:0] local_bb2_and196_i;

assign local_bb2_and196_i_inputs_ready = rnode_173to174_bb2_add193_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and196_i = (rnode_173to174_bb2_add193_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb2_and196_i_valid_out = 1'b1;
assign rnode_173to174_bb2_add193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and199_i_valid_out;
wire local_bb2_and199_i_stall_in;
wire local_bb2_and199_i_inputs_ready;
wire local_bb2_and199_i_stall_local;
wire [31:0] local_bb2_and199_i;

assign local_bb2_and199_i_inputs_ready = rnode_173to174_bb2_add193_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb2_and199_i = (rnode_173to174_bb2_add193_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb2_and199_i_valid_out = 1'b1;
assign rnode_173to174_bb2_add193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and202_i_stall_local;
wire [31:0] local_bb2_and202_i;

assign local_bb2_and202_i = (rnode_173to174_bb2_add193_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_var__u107_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u107_0_stall_in_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u107_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u107_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u107_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u107_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u107_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u107_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_var__u107_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_var__u107_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_var__u107_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_var__u107_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_var__u107_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2_var__u107_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2_var__u107_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_var__u107_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_var__u107_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_174to175_bb2_var__u107_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_var__u107_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_var__u107_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_var__u107_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_var__u107_0_NO_SHIFT_REG = rnode_174to175_bb2_var__u107_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_var__u107_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_var__u107_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2__26_i1679_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1679_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2__26_i1679_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2__26_i1679_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2__26_i1679_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2__26_i1679_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2__26_i1679_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2__26_i1679_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2__26_i1679_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2__26_i1679_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2__26_i1679_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2__26_i1679_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2__26_i1679_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2__26_i1679_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__26_i1679_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1679_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1679_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i1679_0_NO_SHIFT_REG = rnode_175to176_bb2__26_i1679_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2__26_i1679_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i1679_1_NO_SHIFT_REG = rnode_175to176_bb2__26_i1679_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2__26_i1679_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i1679_2_NO_SHIFT_REG = rnode_175to176_bb2__26_i1679_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and194_i1744_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and194_i1744_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and194_i1744_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and194_i1744_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and194_i1744_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i1744_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and194_i1744_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and194_i1744_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and194_i1744_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and194_i1744_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and194_i1744_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and194_i1744),
	.data_out(rnode_174to175_bb2_and194_i1744_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and194_i1744_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and194_i1744_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and194_i1744_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and194_i1744_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and194_i1744_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and194_i1744_stall_in = 1'b0;
assign rnode_174to175_bb2_and194_i1744_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and194_i1744_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and194_i1744_0_NO_SHIFT_REG = rnode_174to175_bb2_and194_i1744_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and194_i1744_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and194_i1744_1_NO_SHIFT_REG = rnode_174to175_bb2_and194_i1744_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and194_i1744_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and194_i1744_2_NO_SHIFT_REG = rnode_174to175_bb2_and194_i1744_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and196_i1745_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i1745_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and196_i1745_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i1745_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and196_i1745_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i1745_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i1745_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i1745_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and196_i1745_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and196_i1745_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and196_i1745_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and196_i1745_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and196_i1745_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and196_i1745),
	.data_out(rnode_174to175_bb2_and196_i1745_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and196_i1745_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and196_i1745_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and196_i1745_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and196_i1745_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and196_i1745_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and196_i1745_stall_in = 1'b0;
assign rnode_174to175_bb2_and196_i1745_0_NO_SHIFT_REG = rnode_174to175_bb2_and196_i1745_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and196_i1745_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and196_i1745_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and199_i1746_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i1746_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and199_i1746_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i1746_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and199_i1746_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i1746_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i1746_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i1746_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and199_i1746_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and199_i1746_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and199_i1746_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and199_i1746_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and199_i1746_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and199_i1746),
	.data_out(rnode_174to175_bb2_and199_i1746_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and199_i1746_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and199_i1746_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and199_i1746_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and199_i1746_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and199_i1746_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and199_i1746_stall_in = 1'b0;
assign rnode_174to175_bb2_and199_i1746_0_NO_SHIFT_REG = rnode_174to175_bb2_and199_i1746_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and199_i1746_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and199_i1746_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i1748_stall_local;
wire [31:0] local_bb2_shr_i_i1748;

assign local_bb2_shr_i_i1748 = (local_bb2_and202_i1747 >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_var__u102_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u102_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u102_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u102_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u102_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u102_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u102_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u102_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_var__u102_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_var__u102_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_var__u102_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_var__u102_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_var__u102_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2_var__u102_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2_var__u102_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_var__u102_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_var__u102_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_var__u102_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_var__u102_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_var__u102_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_var__u102_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u102_0_NO_SHIFT_REG = rnode_175to176_bb2_var__u102_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_var__u102_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u102_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_not_cmp37_i1223_stall_local;
wire local_bb2_not_cmp37_i1223;

assign local_bb2_not_cmp37_i1223 = (rnode_173to175_bb2_cmp37_i1117_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2__26_i1130_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1130_0_stall_in_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1130_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1130_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1130_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1130_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1130_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i1130_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2__26_i1130_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2__26_i1130_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2__26_i1130_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2__26_i1130_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2__26_i1130_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2__26_i1130_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2__26_i1130_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2__26_i1130_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2__26_i1130_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_174to175_bb2__26_i1130_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2__26_i1130_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2__26_i1130_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2__26_i1130_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__26_i1130_0_NO_SHIFT_REG = rnode_174to175_bb2__26_i1130_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__26_i1130_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__26_i1130_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and193_i1195_valid_out;
wire local_bb2_and193_i1195_stall_in;
wire local_bb2_and193_i1195_inputs_ready;
wire local_bb2_and193_i1195_stall_local;
wire [31:0] local_bb2_and193_i1195;

assign local_bb2_and193_i1195_inputs_ready = rnode_173to174_bb2_add192_i1194_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_and193_i1195 = (rnode_173to174_bb2_add192_i1194_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb2_and193_i1195_valid_out = 1'b1;
assign rnode_173to174_bb2_add192_i1194_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and195_i1196_valid_out;
wire local_bb2_and195_i1196_stall_in;
wire local_bb2_and195_i1196_inputs_ready;
wire local_bb2_and195_i1196_stall_local;
wire [31:0] local_bb2_and195_i1196;

assign local_bb2_and195_i1196_inputs_ready = rnode_173to174_bb2_add192_i1194_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and195_i1196 = (rnode_173to174_bb2_add192_i1194_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb2_and195_i1196_valid_out = 1'b1;
assign rnode_173to174_bb2_add192_i1194_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and198_i1197_valid_out;
wire local_bb2_and198_i1197_stall_in;
wire local_bb2_and198_i1197_inputs_ready;
wire local_bb2_and198_i1197_stall_local;
wire [31:0] local_bb2_and198_i1197;

assign local_bb2_and198_i1197_inputs_ready = rnode_173to174_bb2_add192_i1194_0_valid_out_2_NO_SHIFT_REG;
assign local_bb2_and198_i1197 = (rnode_173to174_bb2_add192_i1194_2_NO_SHIFT_REG & 32'h1);
assign local_bb2_and198_i1197_valid_out = 1'b1;
assign rnode_173to174_bb2_add192_i1194_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and201_i1198_stall_local;
wire [31:0] local_bb2_and201_i1198;

assign local_bb2_and201_i1198 = (rnode_173to174_bb2_add192_i1194_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_var__u111_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u111_0_stall_in_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u111_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u111_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u111_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u111_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u111_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u111_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_var__u111_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_var__u111_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_var__u111_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_var__u111_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_var__u111_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2_var__u111_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2_var__u111_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_var__u111_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_var__u111_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_174to175_bb2_var__u111_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_var__u111_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_var__u111_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_var__u111_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_var__u111_0_NO_SHIFT_REG = rnode_174to175_bb2_var__u111_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_var__u111_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_var__u111_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_not_cmp37_i211_stall_local;
wire local_bb2_not_cmp37_i211;

assign local_bb2_not_cmp37_i211 = (rnode_173to175_bb2_cmp37_i105_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2__26_i118_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i118_0_stall_in_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i118_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i118_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i118_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i118_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i118_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__26_i118_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2__26_i118_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2__26_i118_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2__26_i118_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2__26_i118_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2__26_i118_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2__26_i118_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2__26_i118_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2__26_i118_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2__26_i118_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_174to175_bb2__26_i118_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2__26_i118_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2__26_i118_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2__26_i118_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__26_i118_0_NO_SHIFT_REG = rnode_174to175_bb2__26_i118_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__26_i118_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__26_i118_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and193_i183_valid_out;
wire local_bb2_and193_i183_stall_in;
wire local_bb2_and193_i183_inputs_ready;
wire local_bb2_and193_i183_stall_local;
wire [31:0] local_bb2_and193_i183;

assign local_bb2_and193_i183_inputs_ready = rnode_173to174_bb2_add192_i182_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_and193_i183 = (rnode_173to174_bb2_add192_i182_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb2_and193_i183_valid_out = 1'b1;
assign rnode_173to174_bb2_add192_i182_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and195_i184_valid_out;
wire local_bb2_and195_i184_stall_in;
wire local_bb2_and195_i184_inputs_ready;
wire local_bb2_and195_i184_stall_local;
wire [31:0] local_bb2_and195_i184;

assign local_bb2_and195_i184_inputs_ready = rnode_173to174_bb2_add192_i182_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and195_i184 = (rnode_173to174_bb2_add192_i182_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb2_and195_i184_valid_out = 1'b1;
assign rnode_173to174_bb2_add192_i182_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and198_i185_valid_out;
wire local_bb2_and198_i185_stall_in;
wire local_bb2_and198_i185_inputs_ready;
wire local_bb2_and198_i185_stall_local;
wire [31:0] local_bb2_and198_i185;

assign local_bb2_and198_i185_inputs_ready = rnode_173to174_bb2_add192_i182_0_valid_out_2_NO_SHIFT_REG;
assign local_bb2_and198_i185 = (rnode_173to174_bb2_add192_i182_2_NO_SHIFT_REG & 32'h1);
assign local_bb2_and198_i185_valid_out = 1'b1;
assign rnode_173to174_bb2_add192_i182_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and201_i186_stall_local;
wire [31:0] local_bb2_and201_i186;

assign local_bb2_and201_i186 = (rnode_173to174_bb2_add192_i182_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_var__u114_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u114_0_stall_in_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u114_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u114_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u114_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u114_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u114_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_var__u114_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_var__u114_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_var__u114_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_var__u114_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_var__u114_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_var__u114_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(rnode_173to174_bb2_var__u114_0_NO_SHIFT_REG),
	.data_out(rnode_174to175_bb2_var__u114_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_var__u114_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_var__u114_0_reg_175_fifo.DATA_WIDTH = 1;
defparam rnode_174to175_bb2_var__u114_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_var__u114_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_var__u114_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_173to174_bb2_var__u114_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_var__u114_0_NO_SHIFT_REG = rnode_174to175_bb2_var__u114_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_var__u114_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_var__u114_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2__26_i665_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i665_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2__26_i665_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2__26_i665_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2__26_i665_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2__26_i665_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2__26_i665_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2__26_i665_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2__26_i665_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2__26_i665_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2__26_i665_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2__26_i665_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2__26_i665_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2__26_i665_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__26_i665_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i665_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i665_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i665_0_NO_SHIFT_REG = rnode_175to176_bb2__26_i665_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2__26_i665_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i665_1_NO_SHIFT_REG = rnode_175to176_bb2__26_i665_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2__26_i665_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i665_2_NO_SHIFT_REG = rnode_175to176_bb2__26_i665_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and194_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and194_i_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and194_i_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and194_i_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and194_i_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and194_i_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and194_i_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and194_i_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and194_i_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and194_i_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and194_i_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and194_i),
	.data_out(rnode_174to175_bb2_and194_i_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and194_i_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and194_i_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and194_i_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and194_i_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and194_i_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and194_i_stall_in = 1'b0;
assign rnode_174to175_bb2_and194_i_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and194_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and194_i_0_NO_SHIFT_REG = rnode_174to175_bb2_and194_i_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and194_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and194_i_1_NO_SHIFT_REG = rnode_174to175_bb2_and194_i_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and194_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and194_i_2_NO_SHIFT_REG = rnode_174to175_bb2_and194_i_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and196_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and196_i_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and196_i_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and196_i_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and196_i_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and196_i_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and196_i_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and196_i_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and196_i_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and196_i),
	.data_out(rnode_174to175_bb2_and196_i_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and196_i_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and196_i_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and196_i_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and196_i_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and196_i_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and196_i_stall_in = 1'b0;
assign rnode_174to175_bb2_and196_i_0_NO_SHIFT_REG = rnode_174to175_bb2_and196_i_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and196_i_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and196_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and199_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and199_i_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and199_i_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and199_i_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and199_i_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and199_i_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and199_i_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and199_i_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and199_i_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and199_i),
	.data_out(rnode_174to175_bb2_and199_i_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and199_i_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and199_i_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and199_i_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and199_i_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and199_i_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and199_i_stall_in = 1'b0;
assign rnode_174to175_bb2_and199_i_0_NO_SHIFT_REG = rnode_174to175_bb2_and199_i_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and199_i_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and199_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i691_stall_local;
wire [31:0] local_bb2_shr_i_i691;

assign local_bb2_shr_i_i691 = (local_bb2_and202_i >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_var__u107_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u107_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u107_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u107_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u107_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u107_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u107_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u107_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_var__u107_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_var__u107_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_var__u107_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_var__u107_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_var__u107_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2_var__u107_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2_var__u107_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_var__u107_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_var__u107_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_var__u107_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_var__u107_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_var__u107_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_var__u107_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u107_0_NO_SHIFT_REG = rnode_175to176_bb2_var__u107_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_var__u107_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u107_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cond293_i1806_stall_local;
wire [31:0] local_bb2_cond293_i1806;

assign local_bb2_cond293_i1806 = (rnode_175to176_bb2__26_i1679_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u124_stall_local;
wire [31:0] local_bb2_var__u124;

assign local_bb2_var__u124[31:1] = 31'h0;
assign local_bb2_var__u124[0] = rnode_175to176_bb2__26_i1679_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr217_i1769_stall_local;
wire [31:0] local_bb2_shr217_i1769;

assign local_bb2_shr217_i1769 = (rnode_174to175_bb2_and194_i1744_1_NO_SHIFT_REG >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__pre_i1767_stall_local;
wire [31:0] local_bb2__pre_i1767;

assign local_bb2__pre_i1767 = (rnode_174to175_bb2_and196_i1745_0_NO_SHIFT_REG & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i1749_stall_local;
wire [31:0] local_bb2_or_i_i1749;

assign local_bb2_or_i_i1749 = (local_bb2_shr_i_i1748 | local_bb2_and202_i1747);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2__26_i1130_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i1130_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2__26_i1130_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2__26_i1130_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2__26_i1130_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2__26_i1130_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2__26_i1130_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2__26_i1130_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2__26_i1130_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2__26_i1130_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2__26_i1130_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2__26_i1130_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2__26_i1130_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2__26_i1130_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__26_i1130_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1130_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1130_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i1130_0_NO_SHIFT_REG = rnode_175to176_bb2__26_i1130_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2__26_i1130_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i1130_1_NO_SHIFT_REG = rnode_175to176_bb2__26_i1130_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2__26_i1130_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i1130_2_NO_SHIFT_REG = rnode_175to176_bb2__26_i1130_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and193_i1195_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and193_i1195_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and193_i1195_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and193_i1195_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and193_i1195_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i1195_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and193_i1195_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and193_i1195_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and193_i1195_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and193_i1195_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and193_i1195_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and193_i1195),
	.data_out(rnode_174to175_bb2_and193_i1195_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and193_i1195_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and193_i1195_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and193_i1195_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and193_i1195_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and193_i1195_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and193_i1195_stall_in = 1'b0;
assign rnode_174to175_bb2_and193_i1195_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and193_i1195_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and193_i1195_0_NO_SHIFT_REG = rnode_174to175_bb2_and193_i1195_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and193_i1195_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and193_i1195_1_NO_SHIFT_REG = rnode_174to175_bb2_and193_i1195_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and193_i1195_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and193_i1195_2_NO_SHIFT_REG = rnode_174to175_bb2_and193_i1195_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and195_i1196_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i1196_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and195_i1196_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i1196_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and195_i1196_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i1196_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i1196_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i1196_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and195_i1196_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and195_i1196_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and195_i1196_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and195_i1196_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and195_i1196_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and195_i1196),
	.data_out(rnode_174to175_bb2_and195_i1196_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and195_i1196_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and195_i1196_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and195_i1196_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and195_i1196_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and195_i1196_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and195_i1196_stall_in = 1'b0;
assign rnode_174to175_bb2_and195_i1196_0_NO_SHIFT_REG = rnode_174to175_bb2_and195_i1196_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and195_i1196_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and195_i1196_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and198_i1197_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i1197_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and198_i1197_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i1197_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and198_i1197_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i1197_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i1197_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i1197_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and198_i1197_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and198_i1197_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and198_i1197_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and198_i1197_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and198_i1197_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and198_i1197),
	.data_out(rnode_174to175_bb2_and198_i1197_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and198_i1197_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and198_i1197_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and198_i1197_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and198_i1197_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and198_i1197_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and198_i1197_stall_in = 1'b0;
assign rnode_174to175_bb2_and198_i1197_0_NO_SHIFT_REG = rnode_174to175_bb2_and198_i1197_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and198_i1197_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and198_i1197_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i1199_stall_local;
wire [31:0] local_bb2_shr_i_i1199;

assign local_bb2_shr_i_i1199 = (local_bb2_and201_i1198 >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_var__u111_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u111_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u111_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u111_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u111_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u111_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u111_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u111_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_var__u111_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_var__u111_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_var__u111_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_var__u111_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_var__u111_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2_var__u111_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2_var__u111_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_var__u111_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_var__u111_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_var__u111_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_var__u111_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_var__u111_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_var__u111_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u111_0_NO_SHIFT_REG = rnode_175to176_bb2_var__u111_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_var__u111_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u111_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2__26_i118_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_2_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2__26_i118_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2__26_i118_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2__26_i118_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2__26_i118_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2__26_i118_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2__26_i118_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2__26_i118_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2__26_i118_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2__26_i118_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2__26_i118_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2__26_i118_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2__26_i118_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2__26_i118_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__26_i118_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i118_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i118_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i118_0_NO_SHIFT_REG = rnode_175to176_bb2__26_i118_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2__26_i118_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i118_1_NO_SHIFT_REG = rnode_175to176_bb2__26_i118_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2__26_i118_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2__26_i118_2_NO_SHIFT_REG = rnode_175to176_bb2__26_i118_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and193_i183_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and193_i183_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and193_i183_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and193_i183_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and193_i183_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and193_i183_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and193_i183_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and193_i183_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and193_i183_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and193_i183_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and193_i183_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and193_i183),
	.data_out(rnode_174to175_bb2_and193_i183_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and193_i183_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and193_i183_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and193_i183_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and193_i183_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and193_i183_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and193_i183_stall_in = 1'b0;
assign rnode_174to175_bb2_and193_i183_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and193_i183_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and193_i183_0_NO_SHIFT_REG = rnode_174to175_bb2_and193_i183_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and193_i183_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and193_i183_1_NO_SHIFT_REG = rnode_174to175_bb2_and193_i183_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and193_i183_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_and193_i183_2_NO_SHIFT_REG = rnode_174to175_bb2_and193_i183_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and195_i184_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i184_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and195_i184_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i184_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and195_i184_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i184_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i184_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and195_i184_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and195_i184_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and195_i184_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and195_i184_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and195_i184_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and195_i184_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and195_i184),
	.data_out(rnode_174to175_bb2_and195_i184_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and195_i184_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and195_i184_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and195_i184_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and195_i184_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and195_i184_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and195_i184_stall_in = 1'b0;
assign rnode_174to175_bb2_and195_i184_0_NO_SHIFT_REG = rnode_174to175_bb2_and195_i184_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and195_i184_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and195_i184_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2_and198_i185_0_valid_out_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i185_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and198_i185_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i185_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2_and198_i185_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i185_0_valid_out_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i185_0_stall_in_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2_and198_i185_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2_and198_i185_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2_and198_i185_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2_and198_i185_0_stall_in_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2_and198_i185_0_valid_out_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2_and198_i185_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2_and198_i185),
	.data_out(rnode_174to175_bb2_and198_i185_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2_and198_i185_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2_and198_i185_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2_and198_i185_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2_and198_i185_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2_and198_i185_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and198_i185_stall_in = 1'b0;
assign rnode_174to175_bb2_and198_i185_0_NO_SHIFT_REG = rnode_174to175_bb2_and198_i185_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2_and198_i185_0_stall_in_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and198_i185_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i187_stall_local;
wire [31:0] local_bb2_shr_i_i187;

assign local_bb2_shr_i_i187 = (local_bb2_and201_i186 >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_var__u114_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u114_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u114_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u114_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u114_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u114_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u114_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_var__u114_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_var__u114_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_var__u114_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_var__u114_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_var__u114_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_var__u114_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(rnode_174to175_bb2_var__u114_0_NO_SHIFT_REG),
	.data_out(rnode_175to176_bb2_var__u114_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_var__u114_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_var__u114_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_var__u114_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_var__u114_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_var__u114_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2_var__u114_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u114_0_NO_SHIFT_REG = rnode_175to176_bb2_var__u114_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_var__u114_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u114_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cond293_i_stall_local;
wire [31:0] local_bb2_cond293_i;

assign local_bb2_cond293_i = (rnode_175to176_bb2__26_i665_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u125_stall_local;
wire [31:0] local_bb2_var__u125;

assign local_bb2_var__u125[31:1] = 31'h0;
assign local_bb2_var__u125[0] = rnode_175to176_bb2__26_i665_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr217_i_stall_local;
wire [31:0] local_bb2_shr217_i;

assign local_bb2_shr217_i = (rnode_174to175_bb2_and194_i_1_NO_SHIFT_REG >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__pre_i705_stall_local;
wire [31:0] local_bb2__pre_i705;

assign local_bb2__pre_i705 = (rnode_174to175_bb2_and196_i_0_NO_SHIFT_REG & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i692_stall_local;
wire [31:0] local_bb2_or_i_i692;

assign local_bb2_or_i_i692 = (local_bb2_shr_i_i691 | local_bb2_and202_i);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext_i1816_stall_local;
wire [31:0] local_bb2_lnot_ext_i1816;

assign local_bb2_lnot_ext_i1816 = (local_bb2_var__u124 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or220_i1770_stall_local;
wire [31:0] local_bb2_or220_i1770;

assign local_bb2_or220_i1770 = (local_bb2_shr217_i1769 | rnode_174to175_bb2_and199_i1746_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool214_i1768_stall_local;
wire local_bb2_tobool214_i1768;

assign local_bb2_tobool214_i1768 = (local_bb2__pre_i1767 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shr1_i_i1750_stall_local;
wire [31:0] local_bb2_shr1_i_i1750;

assign local_bb2_shr1_i_i1750 = (local_bb2_or_i_i1749 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_cond292_i1257_stall_local;
wire [31:0] local_bb2_cond292_i1257;

assign local_bb2_cond292_i1257 = (rnode_175to176_bb2__26_i1130_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u126_stall_local;
wire [31:0] local_bb2_var__u126;

assign local_bb2_var__u126[31:1] = 31'h0;
assign local_bb2_var__u126[0] = rnode_175to176_bb2__26_i1130_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr216_i1220_stall_local;
wire [31:0] local_bb2_shr216_i1220;

assign local_bb2_shr216_i1220 = (rnode_174to175_bb2_and193_i1195_1_NO_SHIFT_REG >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__pre_i1218_stall_local;
wire [31:0] local_bb2__pre_i1218;

assign local_bb2__pre_i1218 = (rnode_174to175_bb2_and195_i1196_0_NO_SHIFT_REG & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i1200_stall_local;
wire [31:0] local_bb2_or_i_i1200;

assign local_bb2_or_i_i1200 = (local_bb2_shr_i_i1199 | local_bb2_and201_i1198);

// This section implements an unregistered operation.
// 
wire local_bb2_cond292_i245_stall_local;
wire [31:0] local_bb2_cond292_i245;

assign local_bb2_cond292_i245 = (rnode_175to176_bb2__26_i118_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u127_stall_local;
wire [31:0] local_bb2_var__u127;

assign local_bb2_var__u127[31:1] = 31'h0;
assign local_bb2_var__u127[0] = rnode_175to176_bb2__26_i118_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr216_i208_stall_local;
wire [31:0] local_bb2_shr216_i208;

assign local_bb2_shr216_i208 = (rnode_174to175_bb2_and193_i183_1_NO_SHIFT_REG >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__pre_i206_stall_local;
wire [31:0] local_bb2__pre_i206;

assign local_bb2__pre_i206 = (rnode_174to175_bb2_and195_i184_0_NO_SHIFT_REG & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i188_stall_local;
wire [31:0] local_bb2_or_i_i188;

assign local_bb2_or_i_i188 = (local_bb2_shr_i_i187 | local_bb2_and201_i186);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext_i722_stall_local;
wire [31:0] local_bb2_lnot_ext_i722;

assign local_bb2_lnot_ext_i722 = (local_bb2_var__u125 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or220_i_stall_local;
wire [31:0] local_bb2_or220_i;

assign local_bb2_or220_i = (local_bb2_shr217_i | rnode_174to175_bb2_and199_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool214_i_stall_local;
wire local_bb2_tobool214_i;

assign local_bb2_tobool214_i = (local_bb2__pre_i705 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shr1_i_i693_stall_local;
wire [31:0] local_bb2_shr1_i_i693;

assign local_bb2_shr1_i_i693 = (local_bb2_or_i_i692 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2__40_demorgan_i1771_stall_local;
wire local_bb2__40_demorgan_i1771;

assign local_bb2__40_demorgan_i1771 = (rnode_173to175_bb2_cmp38_i1666_0_NO_SHIFT_REG | local_bb2_tobool214_i1768);

// This section implements an unregistered operation.
// 
wire local_bb2__42_i1773_stall_local;
wire local_bb2__42_i1773;

assign local_bb2__42_i1773 = (local_bb2_tobool214_i1768 & local_bb2_not_cmp38_i1772);

// This section implements an unregistered operation.
// 
wire local_bb2_or2_i_i1751_stall_local;
wire [31:0] local_bb2_or2_i_i1751;

assign local_bb2_or2_i_i1751 = (local_bb2_shr1_i_i1750 | local_bb2_or_i_i1749);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext_i1267_stall_local;
wire [31:0] local_bb2_lnot_ext_i1267;

assign local_bb2_lnot_ext_i1267 = (local_bb2_var__u126 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or219_i1221_stall_local;
wire [31:0] local_bb2_or219_i1221;

assign local_bb2_or219_i1221 = (local_bb2_shr216_i1220 | rnode_174to175_bb2_and198_i1197_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool213_i1219_stall_local;
wire local_bb2_tobool213_i1219;

assign local_bb2_tobool213_i1219 = (local_bb2__pre_i1218 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shr1_i_i1201_stall_local;
wire [31:0] local_bb2_shr1_i_i1201;

assign local_bb2_shr1_i_i1201 = (local_bb2_or_i_i1200 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext_i255_stall_local;
wire [31:0] local_bb2_lnot_ext_i255;

assign local_bb2_lnot_ext_i255 = (local_bb2_var__u127 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or219_i209_stall_local;
wire [31:0] local_bb2_or219_i209;

assign local_bb2_or219_i209 = (local_bb2_shr216_i208 | rnode_174to175_bb2_and198_i185_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool213_i207_stall_local;
wire local_bb2_tobool213_i207;

assign local_bb2_tobool213_i207 = (local_bb2__pre_i206 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shr1_i_i189_stall_local;
wire [31:0] local_bb2_shr1_i_i189;

assign local_bb2_shr1_i_i189 = (local_bb2_or_i_i188 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2__40_demorgan_i706_stall_local;
wire local_bb2__40_demorgan_i706;

assign local_bb2__40_demorgan_i706 = (rnode_173to175_bb2_cmp38_i_0_NO_SHIFT_REG | local_bb2_tobool214_i);

// This section implements an unregistered operation.
// 
wire local_bb2__42_i707_stall_local;
wire local_bb2__42_i707;

assign local_bb2__42_i707 = (local_bb2_tobool214_i & local_bb2_not_cmp38_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or2_i_i694_stall_local;
wire [31:0] local_bb2_or2_i_i694;

assign local_bb2_or2_i_i694 = (local_bb2_shr1_i_i693 | local_bb2_or_i_i692);

// This section implements an unregistered operation.
// 
wire local_bb2__43_i1774_stall_local;
wire [31:0] local_bb2__43_i1774;

assign local_bb2__43_i1774 = (local_bb2__42_i1773 ? 32'h0 : local_bb2__pre_i1767);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_i1752_stall_local;
wire [31:0] local_bb2_shr3_i_i1752;

assign local_bb2_shr3_i_i1752 = (local_bb2_or2_i_i1751 >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2__40_demorgan_i1222_stall_local;
wire local_bb2__40_demorgan_i1222;

assign local_bb2__40_demorgan_i1222 = (rnode_173to175_bb2_cmp37_i1117_0_NO_SHIFT_REG | local_bb2_tobool213_i1219);

// This section implements an unregistered operation.
// 
wire local_bb2__42_i1224_stall_local;
wire local_bb2__42_i1224;

assign local_bb2__42_i1224 = (local_bb2_tobool213_i1219 & local_bb2_not_cmp37_i1223);

// This section implements an unregistered operation.
// 
wire local_bb2_or2_i_i1202_stall_local;
wire [31:0] local_bb2_or2_i_i1202;

assign local_bb2_or2_i_i1202 = (local_bb2_shr1_i_i1201 | local_bb2_or_i_i1200);

// This section implements an unregistered operation.
// 
wire local_bb2__40_demorgan_i210_stall_local;
wire local_bb2__40_demorgan_i210;

assign local_bb2__40_demorgan_i210 = (rnode_173to175_bb2_cmp37_i105_0_NO_SHIFT_REG | local_bb2_tobool213_i207);

// This section implements an unregistered operation.
// 
wire local_bb2__42_i212_stall_local;
wire local_bb2__42_i212;

assign local_bb2__42_i212 = (local_bb2_tobool213_i207 & local_bb2_not_cmp37_i211);

// This section implements an unregistered operation.
// 
wire local_bb2_or2_i_i190_stall_local;
wire [31:0] local_bb2_or2_i_i190;

assign local_bb2_or2_i_i190 = (local_bb2_shr1_i_i189 | local_bb2_or_i_i188);

// This section implements an unregistered operation.
// 
wire local_bb2__43_i708_stall_local;
wire [31:0] local_bb2__43_i708;

assign local_bb2__43_i708 = (local_bb2__42_i707 ? 32'h0 : local_bb2__pre_i705);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_i695_stall_local;
wire [31:0] local_bb2_shr3_i_i695;

assign local_bb2_shr3_i_i695 = (local_bb2_or2_i_i694 >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_or4_i_i1753_stall_local;
wire [31:0] local_bb2_or4_i_i1753;

assign local_bb2_or4_i_i1753 = (local_bb2_shr3_i_i1752 | local_bb2_or2_i_i1751);

// This section implements an unregistered operation.
// 
wire local_bb2__43_i1225_stall_local;
wire [31:0] local_bb2__43_i1225;

assign local_bb2__43_i1225 = (local_bb2__42_i1224 ? 32'h0 : local_bb2__pre_i1218);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_i1203_stall_local;
wire [31:0] local_bb2_shr3_i_i1203;

assign local_bb2_shr3_i_i1203 = (local_bb2_or2_i_i1202 >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2__43_i213_stall_local;
wire [31:0] local_bb2__43_i213;

assign local_bb2__43_i213 = (local_bb2__42_i212 ? 32'h0 : local_bb2__pre_i206);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_i191_stall_local;
wire [31:0] local_bb2_shr3_i_i191;

assign local_bb2_shr3_i_i191 = (local_bb2_or2_i_i190 >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_or4_i_i696_stall_local;
wire [31:0] local_bb2_or4_i_i696;

assign local_bb2_or4_i_i696 = (local_bb2_shr3_i_i695 | local_bb2_or2_i_i694);

// This section implements an unregistered operation.
// 
wire local_bb2_shr5_i_i1754_stall_local;
wire [31:0] local_bb2_shr5_i_i1754;

assign local_bb2_shr5_i_i1754 = (local_bb2_or4_i_i1753 >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_or4_i_i1204_stall_local;
wire [31:0] local_bb2_or4_i_i1204;

assign local_bb2_or4_i_i1204 = (local_bb2_shr3_i_i1203 | local_bb2_or2_i_i1202);

// This section implements an unregistered operation.
// 
wire local_bb2_or4_i_i192_stall_local;
wire [31:0] local_bb2_or4_i_i192;

assign local_bb2_or4_i_i192 = (local_bb2_shr3_i_i191 | local_bb2_or2_i_i190);

// This section implements an unregistered operation.
// 
wire local_bb2_shr5_i_i697_stall_local;
wire [31:0] local_bb2_shr5_i_i697;

assign local_bb2_shr5_i_i697 = (local_bb2_or4_i_i696 >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_i_i1755_stall_local;
wire [31:0] local_bb2_or6_i_i1755;

assign local_bb2_or6_i_i1755 = (local_bb2_shr5_i_i1754 | local_bb2_or4_i_i1753);

// This section implements an unregistered operation.
// 
wire local_bb2_shr5_i_i1205_stall_local;
wire [31:0] local_bb2_shr5_i_i1205;

assign local_bb2_shr5_i_i1205 = (local_bb2_or4_i_i1204 >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_shr5_i_i193_stall_local;
wire [31:0] local_bb2_shr5_i_i193;

assign local_bb2_shr5_i_i193 = (local_bb2_or4_i_i192 >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_i_i698_stall_local;
wire [31:0] local_bb2_or6_i_i698;

assign local_bb2_or6_i_i698 = (local_bb2_shr5_i_i697 | local_bb2_or4_i_i696);

// This section implements an unregistered operation.
// 
wire local_bb2_shr7_i_i1756_stall_local;
wire [31:0] local_bb2_shr7_i_i1756;

assign local_bb2_shr7_i_i1756 = (local_bb2_or6_i_i1755 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_masked_i_i1757_stall_local;
wire [31:0] local_bb2_or6_masked_i_i1757;

assign local_bb2_or6_masked_i_i1757 = (local_bb2_or6_i_i1755 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_i_i1206_stall_local;
wire [31:0] local_bb2_or6_i_i1206;

assign local_bb2_or6_i_i1206 = (local_bb2_shr5_i_i1205 | local_bb2_or4_i_i1204);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_i_i194_stall_local;
wire [31:0] local_bb2_or6_i_i194;

assign local_bb2_or6_i_i194 = (local_bb2_shr5_i_i193 | local_bb2_or4_i_i192);

// This section implements an unregistered operation.
// 
wire local_bb2_shr7_i_i699_stall_local;
wire [31:0] local_bb2_shr7_i_i699;

assign local_bb2_shr7_i_i699 = (local_bb2_or6_i_i698 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_masked_i_i700_stall_local;
wire [31:0] local_bb2_or6_masked_i_i700;

assign local_bb2_or6_masked_i_i700 = (local_bb2_or6_i_i698 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_neg_i_i1758_stall_local;
wire [31:0] local_bb2_neg_i_i1758;

assign local_bb2_neg_i_i1758 = (local_bb2_or6_masked_i_i1757 | local_bb2_shr7_i_i1756);

// This section implements an unregistered operation.
// 
wire local_bb2_shr7_i_i1207_stall_local;
wire [31:0] local_bb2_shr7_i_i1207;

assign local_bb2_shr7_i_i1207 = (local_bb2_or6_i_i1206 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_masked_i_i1208_stall_local;
wire [31:0] local_bb2_or6_masked_i_i1208;

assign local_bb2_or6_masked_i_i1208 = (local_bb2_or6_i_i1206 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr7_i_i195_stall_local;
wire [31:0] local_bb2_shr7_i_i195;

assign local_bb2_shr7_i_i195 = (local_bb2_or6_i_i194 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_masked_i_i196_stall_local;
wire [31:0] local_bb2_or6_masked_i_i196;

assign local_bb2_or6_masked_i_i196 = (local_bb2_or6_i_i194 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_neg_i_i701_stall_local;
wire [31:0] local_bb2_neg_i_i701;

assign local_bb2_neg_i_i701 = (local_bb2_or6_masked_i_i700 | local_bb2_shr7_i_i699);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_i1759_stall_local;
wire [31:0] local_bb2_and_i_i1759;

assign local_bb2_and_i_i1759 = (local_bb2_neg_i_i1758 ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_neg_i_i1209_stall_local;
wire [31:0] local_bb2_neg_i_i1209;

assign local_bb2_neg_i_i1209 = (local_bb2_or6_masked_i_i1208 | local_bb2_shr7_i_i1207);

// This section implements an unregistered operation.
// 
wire local_bb2_neg_i_i197_stall_local;
wire [31:0] local_bb2_neg_i_i197;

assign local_bb2_neg_i_i197 = (local_bb2_or6_masked_i_i196 | local_bb2_shr7_i_i195);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_i702_stall_local;
wire [31:0] local_bb2_and_i_i702;

assign local_bb2_and_i_i702 = (local_bb2_neg_i_i701 ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2__and_i_i1759_valid_out;
wire local_bb2__and_i_i1759_stall_in;
wire local_bb2__and_i_i1759_inputs_ready;
wire local_bb2__and_i_i1759_stall_local;
wire [31:0] local_bb2__and_i_i1759;

thirtysix_six_comp local_bb2__and_i_i1759_popcnt_instance (
	.data(local_bb2_and_i_i1759),
	.sum(local_bb2__and_i_i1759)
);


assign local_bb2__and_i_i1759_inputs_ready = rnode_173to174_bb2_add193_i1743_0_valid_out_3_NO_SHIFT_REG;
assign local_bb2__and_i_i1759_valid_out = 1'b1;
assign rnode_173to174_bb2_add193_i1743_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_i1210_stall_local;
wire [31:0] local_bb2_and_i_i1210;

assign local_bb2_and_i_i1210 = (local_bb2_neg_i_i1209 ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_i198_stall_local;
wire [31:0] local_bb2_and_i_i198;

assign local_bb2_and_i_i198 = (local_bb2_neg_i_i197 ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2__and_i_i702_valid_out;
wire local_bb2__and_i_i702_stall_in;
wire local_bb2__and_i_i702_inputs_ready;
wire local_bb2__and_i_i702_stall_local;
wire [31:0] local_bb2__and_i_i702;

thirtysix_six_comp local_bb2__and_i_i702_popcnt_instance (
	.data(local_bb2_and_i_i702),
	.sum(local_bb2__and_i_i702)
);


assign local_bb2__and_i_i702_inputs_ready = rnode_173to174_bb2_add193_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb2__and_i_i702_valid_out = 1'b1;
assign rnode_173to174_bb2_add193_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2__and_i_i1759_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i1759_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i1759_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i1759_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i1759_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1759_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2__and_i_i1759_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2__and_i_i1759_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2__and_i_i1759_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2__and_i_i1759_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2__and_i_i1759_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2__and_i_i1759),
	.data_out(rnode_174to175_bb2__and_i_i1759_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2__and_i_i1759_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2__and_i_i1759_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2__and_i_i1759_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2__and_i_i1759_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2__and_i_i1759_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__and_i_i1759_stall_in = 1'b0;
assign rnode_174to175_bb2__and_i_i1759_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i1759_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i1759_0_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i1759_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__and_i_i1759_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i1759_1_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i1759_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__and_i_i1759_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i1759_2_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i1759_0_reg_175_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__and_i_i1210_valid_out;
wire local_bb2__and_i_i1210_stall_in;
wire local_bb2__and_i_i1210_inputs_ready;
wire local_bb2__and_i_i1210_stall_local;
wire [31:0] local_bb2__and_i_i1210;

thirtysix_six_comp local_bb2__and_i_i1210_popcnt_instance (
	.data(local_bb2_and_i_i1210),
	.sum(local_bb2__and_i_i1210)
);


assign local_bb2__and_i_i1210_inputs_ready = rnode_173to174_bb2_add192_i1194_0_valid_out_3_NO_SHIFT_REG;
assign local_bb2__and_i_i1210_valid_out = 1'b1;
assign rnode_173to174_bb2_add192_i1194_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2__and_i_i198_valid_out;
wire local_bb2__and_i_i198_stall_in;
wire local_bb2__and_i_i198_inputs_ready;
wire local_bb2__and_i_i198_stall_local;
wire [31:0] local_bb2__and_i_i198;

thirtysix_six_comp local_bb2__and_i_i198_popcnt_instance (
	.data(local_bb2_and_i_i198),
	.sum(local_bb2__and_i_i198)
);


assign local_bb2__and_i_i198_inputs_ready = rnode_173to174_bb2_add192_i182_0_valid_out_3_NO_SHIFT_REG;
assign local_bb2__and_i_i198_valid_out = 1'b1;
assign rnode_173to174_bb2_add192_i182_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2__and_i_i702_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i702_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i702_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i702_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i702_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i702_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2__and_i_i702_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2__and_i_i702_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2__and_i_i702_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2__and_i_i702_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2__and_i_i702_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2__and_i_i702),
	.data_out(rnode_174to175_bb2__and_i_i702_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2__and_i_i702_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2__and_i_i702_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2__and_i_i702_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2__and_i_i702_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2__and_i_i702_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__and_i_i702_stall_in = 1'b0;
assign rnode_174to175_bb2__and_i_i702_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i702_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i702_0_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i702_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__and_i_i702_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i702_1_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i702_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__and_i_i702_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i702_2_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i702_0_reg_175_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and9_i_i1760_stall_local;
wire [31:0] local_bb2_and9_i_i1760;

assign local_bb2_and9_i_i1760 = (rnode_174to175_bb2__and_i_i1759_0_NO_SHIFT_REG & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and204_i1761_stall_local;
wire [31:0] local_bb2_and204_i1761;

assign local_bb2_and204_i1761 = (rnode_174to175_bb2__and_i_i1759_1_NO_SHIFT_REG & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_and207_i1763_stall_local;
wire [31:0] local_bb2_and207_i1763;

assign local_bb2_and207_i1763 = (rnode_174to175_bb2__and_i_i1759_2_NO_SHIFT_REG & 32'h7);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2__and_i_i1210_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i1210_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i1210_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i1210_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i1210_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i1210_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2__and_i_i1210_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2__and_i_i1210_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2__and_i_i1210_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2__and_i_i1210_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2__and_i_i1210_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2__and_i_i1210),
	.data_out(rnode_174to175_bb2__and_i_i1210_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2__and_i_i1210_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2__and_i_i1210_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2__and_i_i1210_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2__and_i_i1210_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2__and_i_i1210_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__and_i_i1210_stall_in = 1'b0;
assign rnode_174to175_bb2__and_i_i1210_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i1210_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i1210_0_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i1210_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__and_i_i1210_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i1210_1_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i1210_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__and_i_i1210_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i1210_2_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i1210_0_reg_175_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_174to175_bb2__and_i_i198_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i198_0_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i198_1_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i198_2_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_reg_175_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_174to175_bb2__and_i_i198_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_valid_out_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_stall_in_0_reg_175_NO_SHIFT_REG;
 logic rnode_174to175_bb2__and_i_i198_0_stall_out_reg_175_NO_SHIFT_REG;

acl_data_fifo rnode_174to175_bb2__and_i_i198_0_reg_175_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_174to175_bb2__and_i_i198_0_reg_175_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_174to175_bb2__and_i_i198_0_stall_in_0_reg_175_NO_SHIFT_REG),
	.valid_out(rnode_174to175_bb2__and_i_i198_0_valid_out_0_reg_175_NO_SHIFT_REG),
	.stall_out(rnode_174to175_bb2__and_i_i198_0_stall_out_reg_175_NO_SHIFT_REG),
	.data_in(local_bb2__and_i_i198),
	.data_out(rnode_174to175_bb2__and_i_i198_0_reg_175_NO_SHIFT_REG)
);

defparam rnode_174to175_bb2__and_i_i198_0_reg_175_fifo.DEPTH = 1;
defparam rnode_174to175_bb2__and_i_i198_0_reg_175_fifo.DATA_WIDTH = 32;
defparam rnode_174to175_bb2__and_i_i198_0_reg_175_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_174to175_bb2__and_i_i198_0_reg_175_fifo.IMPL = "shift_reg";

assign rnode_174to175_bb2__and_i_i198_0_reg_175_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__and_i_i198_stall_in = 1'b0;
assign rnode_174to175_bb2__and_i_i198_0_stall_in_0_reg_175_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i198_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i198_0_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i198_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__and_i_i198_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i198_1_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i198_0_reg_175_NO_SHIFT_REG;
assign rnode_174to175_bb2__and_i_i198_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_174to175_bb2__and_i_i198_2_NO_SHIFT_REG = rnode_174to175_bb2__and_i_i198_0_reg_175_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and9_i_i703_stall_local;
wire [31:0] local_bb2_and9_i_i703;

assign local_bb2_and9_i_i703 = (rnode_174to175_bb2__and_i_i702_0_NO_SHIFT_REG & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and204_i_stall_local;
wire [31:0] local_bb2_and204_i;

assign local_bb2_and204_i = (rnode_174to175_bb2__and_i_i702_1_NO_SHIFT_REG & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_and207_i_stall_local;
wire [31:0] local_bb2_and207_i;

assign local_bb2_and207_i = (rnode_174to175_bb2__and_i_i702_2_NO_SHIFT_REG & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_sub240_i1782_stall_local;
wire [31:0] local_bb2_sub240_i1782;

assign local_bb2_sub240_i1782 = (32'h0 - local_bb2_and9_i_i1760);

// This section implements an unregistered operation.
// 
wire local_bb2_shl205_i1762_stall_local;
wire [31:0] local_bb2_shl205_i1762;

assign local_bb2_shl205_i1762 = (rnode_174to175_bb2_and194_i1744_0_NO_SHIFT_REG << local_bb2_and204_i1761);

// This section implements an unregistered operation.
// 
wire local_bb2_and9_i_i1211_stall_local;
wire [31:0] local_bb2_and9_i_i1211;

assign local_bb2_and9_i_i1211 = (rnode_174to175_bb2__and_i_i1210_0_NO_SHIFT_REG & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and203_i1212_stall_local;
wire [31:0] local_bb2_and203_i1212;

assign local_bb2_and203_i1212 = (rnode_174to175_bb2__and_i_i1210_1_NO_SHIFT_REG & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_and206_i1214_stall_local;
wire [31:0] local_bb2_and206_i1214;

assign local_bb2_and206_i1214 = (rnode_174to175_bb2__and_i_i1210_2_NO_SHIFT_REG & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_and9_i_i199_stall_local;
wire [31:0] local_bb2_and9_i_i199;

assign local_bb2_and9_i_i199 = (rnode_174to175_bb2__and_i_i198_0_NO_SHIFT_REG & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and203_i200_stall_local;
wire [31:0] local_bb2_and203_i200;

assign local_bb2_and203_i200 = (rnode_174to175_bb2__and_i_i198_1_NO_SHIFT_REG & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_and206_i202_stall_local;
wire [31:0] local_bb2_and206_i202;

assign local_bb2_and206_i202 = (rnode_174to175_bb2__and_i_i198_2_NO_SHIFT_REG & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_sub240_i_stall_local;
wire [31:0] local_bb2_sub240_i;

assign local_bb2_sub240_i = (32'h0 - local_bb2_and9_i_i703);

// This section implements an unregistered operation.
// 
wire local_bb2_shl205_i_stall_local;
wire [31:0] local_bb2_shl205_i;

assign local_bb2_shl205_i = (rnode_174to175_bb2_and194_i_0_NO_SHIFT_REG << local_bb2_and204_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cond245_i1783_stall_local;
wire [31:0] local_bb2_cond245_i1783;

assign local_bb2_cond245_i1783 = (rnode_173to175_bb2_cmp38_i1666_2_NO_SHIFT_REG ? local_bb2_sub240_i1782 : local_bb2__43_i1774);

// This section implements an unregistered operation.
// 
wire local_bb2_and206_i1764_stall_local;
wire [31:0] local_bb2_and206_i1764;

assign local_bb2_and206_i1764 = (local_bb2_shl205_i1762 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub239_i1233_stall_local;
wire [31:0] local_bb2_sub239_i1233;

assign local_bb2_sub239_i1233 = (32'h0 - local_bb2_and9_i_i1211);

// This section implements an unregistered operation.
// 
wire local_bb2_shl204_i1213_stall_local;
wire [31:0] local_bb2_shl204_i1213;

assign local_bb2_shl204_i1213 = (rnode_174to175_bb2_and193_i1195_0_NO_SHIFT_REG << local_bb2_and203_i1212);

// This section implements an unregistered operation.
// 
wire local_bb2_sub239_i221_stall_local;
wire [31:0] local_bb2_sub239_i221;

assign local_bb2_sub239_i221 = (32'h0 - local_bb2_and9_i_i199);

// This section implements an unregistered operation.
// 
wire local_bb2_shl204_i201_stall_local;
wire [31:0] local_bb2_shl204_i201;

assign local_bb2_shl204_i201 = (rnode_174to175_bb2_and193_i183_0_NO_SHIFT_REG << local_bb2_and203_i200);

// This section implements an unregistered operation.
// 
wire local_bb2_cond245_i_stall_local;
wire [31:0] local_bb2_cond245_i;

assign local_bb2_cond245_i = (rnode_173to175_bb2_cmp38_i_2_NO_SHIFT_REG ? local_bb2_sub240_i : local_bb2__43_i708);

// This section implements an unregistered operation.
// 
wire local_bb2_and206_i704_stall_local;
wire [31:0] local_bb2_and206_i704;

assign local_bb2_and206_i704 = (local_bb2_shl205_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_add246_i1784_stall_local;
wire [31:0] local_bb2_add246_i1784;

assign local_bb2_add246_i1784 = (local_bb2_cond245_i1783 + rnode_173to175_bb2_and17_i1655_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_fold_i1786_stall_local;
wire [31:0] local_bb2_fold_i1786;

assign local_bb2_fold_i1786 = (local_bb2_cond245_i1783 + rnode_173to175_bb2_shr16_i1654_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl208_i1765_stall_local;
wire [31:0] local_bb2_shl208_i1765;

assign local_bb2_shl208_i1765 = (local_bb2_and206_i1764 << local_bb2_and207_i1763);

// This section implements an unregistered operation.
// 
wire local_bb2_cond244_i1234_stall_local;
wire [31:0] local_bb2_cond244_i1234;

assign local_bb2_cond244_i1234 = (rnode_173to175_bb2_cmp37_i1117_2_NO_SHIFT_REG ? local_bb2_sub239_i1233 : local_bb2__43_i1225);

// This section implements an unregistered operation.
// 
wire local_bb2_and205_i1215_stall_local;
wire [31:0] local_bb2_and205_i1215;

assign local_bb2_and205_i1215 = (local_bb2_shl204_i1213 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond244_i222_stall_local;
wire [31:0] local_bb2_cond244_i222;

assign local_bb2_cond244_i222 = (rnode_173to175_bb2_cmp37_i105_2_NO_SHIFT_REG ? local_bb2_sub239_i221 : local_bb2__43_i213);

// This section implements an unregistered operation.
// 
wire local_bb2_and205_i203_stall_local;
wire [31:0] local_bb2_and205_i203;

assign local_bb2_and205_i203 = (local_bb2_shl204_i201 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_add246_i_stall_local;
wire [31:0] local_bb2_add246_i;

assign local_bb2_add246_i = (local_bb2_cond245_i + rnode_173to175_bb2_and17_i643_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_fold_i713_stall_local;
wire [31:0] local_bb2_fold_i713;

assign local_bb2_fold_i713 = (local_bb2_cond245_i + rnode_173to175_bb2_shr16_i642_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl208_i_stall_local;
wire [31:0] local_bb2_shl208_i;

assign local_bb2_shl208_i = (local_bb2_and206_i704 << local_bb2_and207_i);

// This section implements an unregistered operation.
// 
wire local_bb2_and251_i1787_stall_local;
wire [31:0] local_bb2_and251_i1787;

assign local_bb2_and251_i1787 = (local_bb2_fold_i1786 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i1798_stall_local;
wire [31:0] local_bb2_and270_i1798;

assign local_bb2_and270_i1798 = (local_bb2_fold_i1786 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and209_i1766_stall_local;
wire [31:0] local_bb2_and209_i1766;

assign local_bb2_and209_i1766 = (local_bb2_shl208_i1765 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_add245_i1235_stall_local;
wire [31:0] local_bb2_add245_i1235;

assign local_bb2_add245_i1235 = (local_bb2_cond244_i1234 + rnode_173to175_bb2_and17_i1106_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_fold_i1237_stall_local;
wire [31:0] local_bb2_fold_i1237;

assign local_bb2_fold_i1237 = (local_bb2_cond244_i1234 + rnode_173to175_bb2_shr16_i1105_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl207_i1216_stall_local;
wire [31:0] local_bb2_shl207_i1216;

assign local_bb2_shl207_i1216 = (local_bb2_and205_i1215 << local_bb2_and206_i1214);

// This section implements an unregistered operation.
// 
wire local_bb2_add245_i223_stall_local;
wire [31:0] local_bb2_add245_i223;

assign local_bb2_add245_i223 = (local_bb2_cond244_i222 + rnode_173to175_bb2_and17_i94_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_fold_i225_stall_local;
wire [31:0] local_bb2_fold_i225;

assign local_bb2_fold_i225 = (local_bb2_cond244_i222 + rnode_173to175_bb2_shr16_i93_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl207_i204_stall_local;
wire [31:0] local_bb2_shl207_i204;

assign local_bb2_shl207_i204 = (local_bb2_and205_i203 << local_bb2_and206_i202);

// This section implements an unregistered operation.
// 
wire local_bb2_and248_i_stall_local;
wire [31:0] local_bb2_and248_i;

assign local_bb2_and248_i = (local_bb2_add246_i & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb2_and251_i_stall_local;
wire [31:0] local_bb2_and251_i;

assign local_bb2_and251_i = (local_bb2_fold_i713 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i718_stall_local;
wire [31:0] local_bb2_and270_i718;

assign local_bb2_and270_i718 = (local_bb2_fold_i713 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and209_i_stall_local;
wire [31:0] local_bb2_and209_i;

assign local_bb2_and209_i = (local_bb2_shl208_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_notrhs_i1789_stall_local;
wire local_bb2_notrhs_i1789;

assign local_bb2_notrhs_i1789 = (local_bb2_and251_i1787 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__44_i1775_stall_local;
wire [31:0] local_bb2__44_i1775;

assign local_bb2__44_i1775 = (local_bb2__40_demorgan_i1771 ? local_bb2_and209_i1766 : local_bb2_or220_i1770);

// This section implements an unregistered operation.
// 
wire local_bb2_and250_i1238_stall_local;
wire [31:0] local_bb2_and250_i1238;

assign local_bb2_and250_i1238 = (local_bb2_fold_i1237 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i1249_stall_local;
wire [31:0] local_bb2_and269_i1249;

assign local_bb2_and269_i1249 = (local_bb2_fold_i1237 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and208_i1217_stall_local;
wire [31:0] local_bb2_and208_i1217;

assign local_bb2_and208_i1217 = (local_bb2_shl207_i1216 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and250_i226_stall_local;
wire [31:0] local_bb2_and250_i226;

assign local_bb2_and250_i226 = (local_bb2_fold_i225 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i237_stall_local;
wire [31:0] local_bb2_and269_i237;

assign local_bb2_and269_i237 = (local_bb2_fold_i225 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and208_i205_stall_local;
wire [31:0] local_bb2_and208_i205;

assign local_bb2_and208_i205 = (local_bb2_shl207_i204 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_notlhs_i714_stall_local;
wire local_bb2_notlhs_i714;

assign local_bb2_notlhs_i714 = (local_bb2_and248_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_notrhs_i715_stall_local;
wire local_bb2_notrhs_i715;

assign local_bb2_notrhs_i715 = (local_bb2_and251_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__44_i709_stall_local;
wire [31:0] local_bb2__44_i709;

assign local_bb2__44_i709 = (local_bb2__40_demorgan_i706 ? local_bb2_and209_i : local_bb2_or220_i);

// This section implements an unregistered operation.
// 
wire local_bb2__45_i1776_stall_local;
wire [31:0] local_bb2__45_i1776;

assign local_bb2__45_i1776 = (local_bb2__42_i1773 ? rnode_174to175_bb2_and194_i1744_2_NO_SHIFT_REG : local_bb2__44_i1775);

// This section implements an unregistered operation.
// 
wire local_bb2_notrhs_i1240_stall_local;
wire local_bb2_notrhs_i1240;

assign local_bb2_notrhs_i1240 = (local_bb2_and250_i1238 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__44_i1226_stall_local;
wire [31:0] local_bb2__44_i1226;

assign local_bb2__44_i1226 = (local_bb2__40_demorgan_i1222 ? local_bb2_and208_i1217 : local_bb2_or219_i1221);

// This section implements an unregistered operation.
// 
wire local_bb2_notrhs_i228_stall_local;
wire local_bb2_notrhs_i228;

assign local_bb2_notrhs_i228 = (local_bb2_and250_i226 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__44_i214_stall_local;
wire [31:0] local_bb2__44_i214;

assign local_bb2__44_i214 = (local_bb2__40_demorgan_i210 ? local_bb2_and208_i205 : local_bb2_or219_i209);

// This section implements an unregistered operation.
// 
wire local_bb2_not__46_i716_stall_local;
wire local_bb2_not__46_i716;

assign local_bb2_not__46_i716 = (local_bb2_notrhs_i715 | local_bb2_notlhs_i714);

// This section implements an unregistered operation.
// 
wire local_bb2__45_i710_stall_local;
wire [31:0] local_bb2__45_i710;

assign local_bb2__45_i710 = (local_bb2__42_i707 ? rnode_174to175_bb2_and194_i_2_NO_SHIFT_REG : local_bb2__44_i709);

// This section implements an unregistered operation.
// 
wire local_bb2_and226_i1777_stall_local;
wire [31:0] local_bb2_and226_i1777;

assign local_bb2_and226_i1777 = (local_bb2__45_i1776 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and271_i1795_stall_local;
wire [31:0] local_bb2_and271_i1795;

assign local_bb2_and271_i1795 = (local_bb2__45_i1776 & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_shr272_i1796_stall_local;
wire [31:0] local_bb2_shr272_i1796;

assign local_bb2_shr272_i1796 = (local_bb2__45_i1776 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2__45_i1227_stall_local;
wire [31:0] local_bb2__45_i1227;

assign local_bb2__45_i1227 = (local_bb2__42_i1224 ? rnode_174to175_bb2_and193_i1195_2_NO_SHIFT_REG : local_bb2__44_i1226);

// This section implements an unregistered operation.
// 
wire local_bb2__45_i215_stall_local;
wire [31:0] local_bb2__45_i215;

assign local_bb2__45_i215 = (local_bb2__42_i212 ? rnode_174to175_bb2_and193_i183_2_NO_SHIFT_REG : local_bb2__44_i214);

// This section implements an unregistered operation.
// 
wire local_bb2_and226_i_stall_local;
wire [31:0] local_bb2_and226_i;

assign local_bb2_and226_i = (local_bb2__45_i710 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and271_i_stall_local;
wire [31:0] local_bb2_and271_i;

assign local_bb2_and271_i = (local_bb2__45_i710 & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_shr272_i_stall_local;
wire [31:0] local_bb2_shr272_i;

assign local_bb2_shr272_i = (local_bb2__45_i710 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp227_i1778_stall_local;
wire local_bb2_cmp227_i1778;

assign local_bb2_cmp227_i1778 = (local_bb2_and226_i1777 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp297_i1810_stall_local;
wire local_bb2_cmp297_i1810;

assign local_bb2_cmp297_i1810 = (local_bb2_and271_i1795 > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i1798_valid_out;
wire local_bb2_and270_i1798_stall_in;
 reg local_bb2_and270_i1798_consumed_0_NO_SHIFT_REG;
wire local_bb2_add246_i1784_valid_out;
wire local_bb2_add246_i1784_stall_in;
 reg local_bb2_add246_i1784_consumed_0_NO_SHIFT_REG;
wire local_bb2_notrhs_i1789_valid_out;
wire local_bb2_notrhs_i1789_stall_in;
 reg local_bb2_notrhs_i1789_consumed_0_NO_SHIFT_REG;
wire local_bb2_not_cmp38_i1772_valid_out_1;
wire local_bb2_not_cmp38_i1772_stall_in_1;
 reg local_bb2_not_cmp38_i1772_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr272_i1796_valid_out;
wire local_bb2_shr272_i1796_stall_in;
 reg local_bb2_shr272_i1796_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp227_i1778_valid_out;
wire local_bb2_cmp227_i1778_stall_in;
 reg local_bb2_cmp227_i1778_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp297_i1810_valid_out;
wire local_bb2_cmp297_i1810_stall_in;
 reg local_bb2_cmp297_i1810_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp300_i1811_valid_out;
wire local_bb2_cmp300_i1811_stall_in;
 reg local_bb2_cmp300_i1811_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp300_i1811_inputs_ready;
wire local_bb2_cmp300_i1811_stall_local;
wire local_bb2_cmp300_i1811;

assign local_bb2_cmp300_i1811_inputs_ready = (rnode_173to175_bb2_shr16_i1654_0_valid_out_NO_SHIFT_REG & rnode_173to175_bb2_cmp38_i1666_0_valid_out_2_NO_SHIFT_REG & rnode_173to175_bb2_and17_i1655_0_valid_out_NO_SHIFT_REG & rnode_173to175_bb2_cmp38_i1666_0_valid_out_0_NO_SHIFT_REG & rnode_174to175_bb2_and194_i1744_0_valid_out_2_NO_SHIFT_REG & rnode_173to175_bb2_cmp38_i1666_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2_and196_i1745_0_valid_out_NO_SHIFT_REG & rnode_174to175_bb2_and194_i1744_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2_and199_i1746_0_valid_out_NO_SHIFT_REG & rnode_174to175_bb2_and194_i1744_0_valid_out_0_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i1759_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i1759_0_valid_out_2_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i1759_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_cmp300_i1811 = (local_bb2_and271_i1795 == 32'h4);
assign local_bb2_and270_i1798_valid_out = 1'b1;
assign local_bb2_add246_i1784_valid_out = 1'b1;
assign local_bb2_notrhs_i1789_valid_out = 1'b1;
assign local_bb2_not_cmp38_i1772_valid_out_1 = 1'b1;
assign local_bb2_shr272_i1796_valid_out = 1'b1;
assign local_bb2_cmp227_i1778_valid_out = 1'b1;
assign local_bb2_cmp297_i1810_valid_out = 1'b1;
assign local_bb2_cmp300_i1811_valid_out = 1'b1;
assign rnode_173to175_bb2_shr16_i1654_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp38_i1666_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_and17_i1655_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp38_i1666_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and194_i1744_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp38_i1666_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and196_i1745_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and194_i1744_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and199_i1746_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and194_i1744_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i1759_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i1759_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i1759_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_and270_i1798_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add246_i1784_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_notrhs_i1789_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_not_cmp38_i1772_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr272_i1796_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp227_i1778_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp297_i1810_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp300_i1811_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_and270_i1798_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i1811_inputs_ready & (local_bb2_and270_i1798_consumed_0_NO_SHIFT_REG | ~(local_bb2_and270_i1798_stall_in)) & local_bb2_cmp300_i1811_stall_local);
		local_bb2_add246_i1784_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i1811_inputs_ready & (local_bb2_add246_i1784_consumed_0_NO_SHIFT_REG | ~(local_bb2_add246_i1784_stall_in)) & local_bb2_cmp300_i1811_stall_local);
		local_bb2_notrhs_i1789_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i1811_inputs_ready & (local_bb2_notrhs_i1789_consumed_0_NO_SHIFT_REG | ~(local_bb2_notrhs_i1789_stall_in)) & local_bb2_cmp300_i1811_stall_local);
		local_bb2_not_cmp38_i1772_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp300_i1811_inputs_ready & (local_bb2_not_cmp38_i1772_consumed_1_NO_SHIFT_REG | ~(local_bb2_not_cmp38_i1772_stall_in_1)) & local_bb2_cmp300_i1811_stall_local);
		local_bb2_shr272_i1796_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i1811_inputs_ready & (local_bb2_shr272_i1796_consumed_0_NO_SHIFT_REG | ~(local_bb2_shr272_i1796_stall_in)) & local_bb2_cmp300_i1811_stall_local);
		local_bb2_cmp227_i1778_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i1811_inputs_ready & (local_bb2_cmp227_i1778_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp227_i1778_stall_in)) & local_bb2_cmp300_i1811_stall_local);
		local_bb2_cmp297_i1810_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i1811_inputs_ready & (local_bb2_cmp297_i1810_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp297_i1810_stall_in)) & local_bb2_cmp300_i1811_stall_local);
		local_bb2_cmp300_i1811_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i1811_inputs_ready & (local_bb2_cmp300_i1811_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp300_i1811_stall_in)) & local_bb2_cmp300_i1811_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_and225_i1228_stall_local;
wire [31:0] local_bb2_and225_i1228;

assign local_bb2_and225_i1228 = (local_bb2__45_i1227 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i1246_stall_local;
wire [31:0] local_bb2_and270_i1246;

assign local_bb2_and270_i1246 = (local_bb2__45_i1227 & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_shr271_i1247_stall_local;
wire [31:0] local_bb2_shr271_i1247;

assign local_bb2_shr271_i1247 = (local_bb2__45_i1227 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and225_i216_stall_local;
wire [31:0] local_bb2_and225_i216;

assign local_bb2_and225_i216 = (local_bb2__45_i215 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i234_stall_local;
wire [31:0] local_bb2_and270_i234;

assign local_bb2_and270_i234 = (local_bb2__45_i215 & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_shr271_i235_stall_local;
wire [31:0] local_bb2_shr271_i235;

assign local_bb2_shr271_i235 = (local_bb2__45_i215 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp227_i_stall_local;
wire local_bb2_cmp227_i;

assign local_bb2_cmp227_i = (local_bb2_and226_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp297_i_stall_local;
wire local_bb2_cmp297_i;

assign local_bb2_cmp297_i = (local_bb2_and271_i > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i718_valid_out;
wire local_bb2_and270_i718_stall_in;
 reg local_bb2_and270_i718_consumed_0_NO_SHIFT_REG;
wire local_bb2_add246_i_valid_out_1;
wire local_bb2_add246_i_stall_in_1;
 reg local_bb2_add246_i_consumed_1_NO_SHIFT_REG;
wire local_bb2_not__46_i716_valid_out;
wire local_bb2_not__46_i716_stall_in;
 reg local_bb2_not__46_i716_consumed_0_NO_SHIFT_REG;
wire local_bb2_not_cmp38_i_valid_out_1;
wire local_bb2_not_cmp38_i_stall_in_1;
 reg local_bb2_not_cmp38_i_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr272_i_valid_out;
wire local_bb2_shr272_i_stall_in;
 reg local_bb2_shr272_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp227_i_valid_out;
wire local_bb2_cmp227_i_stall_in;
 reg local_bb2_cmp227_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp297_i_valid_out;
wire local_bb2_cmp297_i_stall_in;
 reg local_bb2_cmp297_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp300_i_valid_out;
wire local_bb2_cmp300_i_stall_in;
 reg local_bb2_cmp300_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp300_i_inputs_ready;
wire local_bb2_cmp300_i_stall_local;
wire local_bb2_cmp300_i;

assign local_bb2_cmp300_i_inputs_ready = (rnode_173to175_bb2_shr16_i642_0_valid_out_NO_SHIFT_REG & rnode_173to175_bb2_cmp38_i_0_valid_out_2_NO_SHIFT_REG & rnode_173to175_bb2_and17_i643_0_valid_out_NO_SHIFT_REG & rnode_173to175_bb2_cmp38_i_0_valid_out_0_NO_SHIFT_REG & rnode_174to175_bb2_and194_i_0_valid_out_2_NO_SHIFT_REG & rnode_173to175_bb2_cmp38_i_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2_and196_i_0_valid_out_NO_SHIFT_REG & rnode_174to175_bb2_and194_i_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2_and199_i_0_valid_out_NO_SHIFT_REG & rnode_174to175_bb2_and194_i_0_valid_out_0_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i702_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i702_0_valid_out_2_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i702_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_cmp300_i = (local_bb2_and271_i == 32'h4);
assign local_bb2_and270_i718_valid_out = 1'b1;
assign local_bb2_add246_i_valid_out_1 = 1'b1;
assign local_bb2_not__46_i716_valid_out = 1'b1;
assign local_bb2_not_cmp38_i_valid_out_1 = 1'b1;
assign local_bb2_shr272_i_valid_out = 1'b1;
assign local_bb2_cmp227_i_valid_out = 1'b1;
assign local_bb2_cmp297_i_valid_out = 1'b1;
assign local_bb2_cmp300_i_valid_out = 1'b1;
assign rnode_173to175_bb2_shr16_i642_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp38_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_and17_i643_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp38_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and194_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp38_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and196_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and194_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and199_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and194_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i702_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i702_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i702_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_and270_i718_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add246_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_not__46_i716_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_not_cmp38_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr272_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp227_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp297_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp300_i_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_and270_i718_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i_inputs_ready & (local_bb2_and270_i718_consumed_0_NO_SHIFT_REG | ~(local_bb2_and270_i718_stall_in)) & local_bb2_cmp300_i_stall_local);
		local_bb2_add246_i_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp300_i_inputs_ready & (local_bb2_add246_i_consumed_1_NO_SHIFT_REG | ~(local_bb2_add246_i_stall_in_1)) & local_bb2_cmp300_i_stall_local);
		local_bb2_not__46_i716_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i_inputs_ready & (local_bb2_not__46_i716_consumed_0_NO_SHIFT_REG | ~(local_bb2_not__46_i716_stall_in)) & local_bb2_cmp300_i_stall_local);
		local_bb2_not_cmp38_i_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp300_i_inputs_ready & (local_bb2_not_cmp38_i_consumed_1_NO_SHIFT_REG | ~(local_bb2_not_cmp38_i_stall_in_1)) & local_bb2_cmp300_i_stall_local);
		local_bb2_shr272_i_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i_inputs_ready & (local_bb2_shr272_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_shr272_i_stall_in)) & local_bb2_cmp300_i_stall_local);
		local_bb2_cmp227_i_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i_inputs_ready & (local_bb2_cmp227_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp227_i_stall_in)) & local_bb2_cmp300_i_stall_local);
		local_bb2_cmp297_i_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i_inputs_ready & (local_bb2_cmp297_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp297_i_stall_in)) & local_bb2_cmp300_i_stall_local);
		local_bb2_cmp300_i_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp300_i_inputs_ready & (local_bb2_cmp300_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp300_i_stall_in)) & local_bb2_cmp300_i_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_and270_i1798_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i1798_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and270_i1798_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i1798_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and270_i1798_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i1798_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i1798_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i1798_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_and270_i1798_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_and270_i1798_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_and270_i1798_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_and270_i1798_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_and270_i1798_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_and270_i1798),
	.data_out(rnode_175to176_bb2_and270_i1798_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_and270_i1798_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_and270_i1798_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_and270_i1798_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_and270_i1798_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_and270_i1798_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and270_i1798_stall_in = 1'b0;
assign rnode_175to176_bb2_and270_i1798_0_NO_SHIFT_REG = rnode_175to176_bb2_and270_i1798_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_and270_i1798_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and270_i1798_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_add246_i1784_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i1784_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add246_i1784_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i1784_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i1784_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add246_i1784_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i1784_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add246_i1784_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i1784_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i1784_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i1784_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_add246_i1784_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_add246_i1784_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_add246_i1784_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_add246_i1784_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_add246_i1784_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_add246_i1784),
	.data_out(rnode_175to176_bb2_add246_i1784_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_add246_i1784_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_add246_i1784_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_add246_i1784_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_add246_i1784_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_add246_i1784_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add246_i1784_stall_in = 1'b0;
assign rnode_175to176_bb2_add246_i1784_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add246_i1784_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_add246_i1784_0_NO_SHIFT_REG = rnode_175to176_bb2_add246_i1784_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_add246_i1784_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_add246_i1784_1_NO_SHIFT_REG = rnode_175to176_bb2_add246_i1784_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_notrhs_i1789_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1789_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1789_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1789_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1789_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1789_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1789_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1789_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_notrhs_i1789_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_notrhs_i1789_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_notrhs_i1789_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_notrhs_i1789_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_notrhs_i1789_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_notrhs_i1789),
	.data_out(rnode_175to176_bb2_notrhs_i1789_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_notrhs_i1789_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_notrhs_i1789_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_notrhs_i1789_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_notrhs_i1789_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_notrhs_i1789_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_notrhs_i1789_stall_in = 1'b0;
assign rnode_175to176_bb2_notrhs_i1789_0_NO_SHIFT_REG = rnode_175to176_bb2_notrhs_i1789_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_notrhs_i1789_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_notrhs_i1789_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_not_cmp38_i1772_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i1772_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i1772_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i1772_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i1772_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i1772_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_not_cmp38_i1772_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_not_cmp38_i1772_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_not_cmp38_i1772_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_not_cmp38_i1772),
	.data_out(rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not_cmp38_i1772_stall_in_1 = 1'b0;
assign rnode_175to176_bb2_not_cmp38_i1772_0_NO_SHIFT_REG = rnode_175to176_bb2_not_cmp38_i1772_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_not_cmp38_i1772_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not_cmp38_i1772_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_shr272_i1796_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i1796_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_shr272_i1796_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i1796_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_shr272_i1796_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i1796_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i1796_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i1796_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_shr272_i1796_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_shr272_i1796_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_shr272_i1796_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_shr272_i1796_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_shr272_i1796_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_shr272_i1796),
	.data_out(rnode_175to176_bb2_shr272_i1796_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_shr272_i1796_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_shr272_i1796_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_shr272_i1796_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_shr272_i1796_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_shr272_i1796_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr272_i1796_stall_in = 1'b0;
assign rnode_175to176_bb2_shr272_i1796_0_NO_SHIFT_REG = rnode_175to176_bb2_shr272_i1796_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_shr272_i1796_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_shr272_i1796_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp227_i1778_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i1778_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp227_i1778_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp227_i1778_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp227_i1778_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp227_i1778_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp227_i1778_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp227_i1778),
	.data_out(rnode_175to176_bb2_cmp227_i1778_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp227_i1778_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp227_i1778_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp227_i1778_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp227_i1778_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp227_i1778_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp227_i1778_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp227_i1778_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp227_i1778_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_cmp227_i1778_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp227_i1778_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp227_i1778_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_cmp227_i1778_1_NO_SHIFT_REG = rnode_175to176_bb2_cmp227_i1778_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp297_i1810_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i1810_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i1810_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i1810_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i1810_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i1810_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i1810_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i1810_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp297_i1810_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp297_i1810_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp297_i1810_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp297_i1810_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp297_i1810_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp297_i1810),
	.data_out(rnode_175to176_bb2_cmp297_i1810_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp297_i1810_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp297_i1810_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp297_i1810_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp297_i1810_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp297_i1810_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp297_i1810_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp297_i1810_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp297_i1810_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp297_i1810_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp297_i1810_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp300_i1811_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i1811_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i1811_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i1811_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i1811_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i1811_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i1811_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i1811_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp300_i1811_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp300_i1811_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp300_i1811_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp300_i1811_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp300_i1811_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp300_i1811),
	.data_out(rnode_175to176_bb2_cmp300_i1811_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp300_i1811_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp300_i1811_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp300_i1811_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp300_i1811_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp300_i1811_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp300_i1811_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp300_i1811_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp300_i1811_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp300_i1811_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp300_i1811_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_i1229_stall_local;
wire local_bb2_cmp226_i1229;

assign local_bb2_cmp226_i1229 = (local_bb2_and225_i1228 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp296_i1261_stall_local;
wire local_bb2_cmp296_i1261;

assign local_bb2_cmp296_i1261 = (local_bb2_and270_i1246 > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i1249_valid_out;
wire local_bb2_and269_i1249_stall_in;
 reg local_bb2_and269_i1249_consumed_0_NO_SHIFT_REG;
wire local_bb2_add245_i1235_valid_out;
wire local_bb2_add245_i1235_stall_in;
 reg local_bb2_add245_i1235_consumed_0_NO_SHIFT_REG;
wire local_bb2_notrhs_i1240_valid_out;
wire local_bb2_notrhs_i1240_stall_in;
 reg local_bb2_notrhs_i1240_consumed_0_NO_SHIFT_REG;
wire local_bb2_not_cmp37_i1223_valid_out_1;
wire local_bb2_not_cmp37_i1223_stall_in_1;
 reg local_bb2_not_cmp37_i1223_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr271_i1247_valid_out;
wire local_bb2_shr271_i1247_stall_in;
 reg local_bb2_shr271_i1247_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp226_i1229_valid_out;
wire local_bb2_cmp226_i1229_stall_in;
 reg local_bb2_cmp226_i1229_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp296_i1261_valid_out;
wire local_bb2_cmp296_i1261_stall_in;
 reg local_bb2_cmp296_i1261_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i1262_valid_out;
wire local_bb2_cmp299_i1262_stall_in;
 reg local_bb2_cmp299_i1262_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i1262_inputs_ready;
wire local_bb2_cmp299_i1262_stall_local;
wire local_bb2_cmp299_i1262;

assign local_bb2_cmp299_i1262_inputs_ready = (rnode_173to175_bb2_shr16_i1105_0_valid_out_NO_SHIFT_REG & rnode_173to175_bb2_cmp37_i1117_0_valid_out_2_NO_SHIFT_REG & rnode_173to175_bb2_and17_i1106_0_valid_out_NO_SHIFT_REG & rnode_173to175_bb2_cmp37_i1117_0_valid_out_0_NO_SHIFT_REG & rnode_174to175_bb2_and193_i1195_0_valid_out_2_NO_SHIFT_REG & rnode_173to175_bb2_cmp37_i1117_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2_and195_i1196_0_valid_out_NO_SHIFT_REG & rnode_174to175_bb2_and193_i1195_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2_and198_i1197_0_valid_out_NO_SHIFT_REG & rnode_174to175_bb2_and193_i1195_0_valid_out_0_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i1210_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i1210_0_valid_out_2_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i1210_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_cmp299_i1262 = (local_bb2_and270_i1246 == 32'h4);
assign local_bb2_and269_i1249_valid_out = 1'b1;
assign local_bb2_add245_i1235_valid_out = 1'b1;
assign local_bb2_notrhs_i1240_valid_out = 1'b1;
assign local_bb2_not_cmp37_i1223_valid_out_1 = 1'b1;
assign local_bb2_shr271_i1247_valid_out = 1'b1;
assign local_bb2_cmp226_i1229_valid_out = 1'b1;
assign local_bb2_cmp296_i1261_valid_out = 1'b1;
assign local_bb2_cmp299_i1262_valid_out = 1'b1;
assign rnode_173to175_bb2_shr16_i1105_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp37_i1117_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_and17_i1106_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp37_i1117_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and193_i1195_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp37_i1117_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and195_i1196_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and193_i1195_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and198_i1197_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and193_i1195_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i1210_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i1210_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i1210_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_and269_i1249_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add245_i1235_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_notrhs_i1240_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_not_cmp37_i1223_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr271_i1247_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp226_i1229_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp296_i1261_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp299_i1262_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_and269_i1249_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1262_inputs_ready & (local_bb2_and269_i1249_consumed_0_NO_SHIFT_REG | ~(local_bb2_and269_i1249_stall_in)) & local_bb2_cmp299_i1262_stall_local);
		local_bb2_add245_i1235_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1262_inputs_ready & (local_bb2_add245_i1235_consumed_0_NO_SHIFT_REG | ~(local_bb2_add245_i1235_stall_in)) & local_bb2_cmp299_i1262_stall_local);
		local_bb2_notrhs_i1240_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1262_inputs_ready & (local_bb2_notrhs_i1240_consumed_0_NO_SHIFT_REG | ~(local_bb2_notrhs_i1240_stall_in)) & local_bb2_cmp299_i1262_stall_local);
		local_bb2_not_cmp37_i1223_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp299_i1262_inputs_ready & (local_bb2_not_cmp37_i1223_consumed_1_NO_SHIFT_REG | ~(local_bb2_not_cmp37_i1223_stall_in_1)) & local_bb2_cmp299_i1262_stall_local);
		local_bb2_shr271_i1247_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1262_inputs_ready & (local_bb2_shr271_i1247_consumed_0_NO_SHIFT_REG | ~(local_bb2_shr271_i1247_stall_in)) & local_bb2_cmp299_i1262_stall_local);
		local_bb2_cmp226_i1229_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1262_inputs_ready & (local_bb2_cmp226_i1229_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp226_i1229_stall_in)) & local_bb2_cmp299_i1262_stall_local);
		local_bb2_cmp296_i1261_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1262_inputs_ready & (local_bb2_cmp296_i1261_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp296_i1261_stall_in)) & local_bb2_cmp299_i1262_stall_local);
		local_bb2_cmp299_i1262_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1262_inputs_ready & (local_bb2_cmp299_i1262_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp299_i1262_stall_in)) & local_bb2_cmp299_i1262_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_i217_stall_local;
wire local_bb2_cmp226_i217;

assign local_bb2_cmp226_i217 = (local_bb2_and225_i216 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp296_i249_stall_local;
wire local_bb2_cmp296_i249;

assign local_bb2_cmp296_i249 = (local_bb2_and270_i234 > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i237_valid_out;
wire local_bb2_and269_i237_stall_in;
 reg local_bb2_and269_i237_consumed_0_NO_SHIFT_REG;
wire local_bb2_add245_i223_valid_out;
wire local_bb2_add245_i223_stall_in;
 reg local_bb2_add245_i223_consumed_0_NO_SHIFT_REG;
wire local_bb2_notrhs_i228_valid_out;
wire local_bb2_notrhs_i228_stall_in;
 reg local_bb2_notrhs_i228_consumed_0_NO_SHIFT_REG;
wire local_bb2_not_cmp37_i211_valid_out_1;
wire local_bb2_not_cmp37_i211_stall_in_1;
 reg local_bb2_not_cmp37_i211_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr271_i235_valid_out;
wire local_bb2_shr271_i235_stall_in;
 reg local_bb2_shr271_i235_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp226_i217_valid_out;
wire local_bb2_cmp226_i217_stall_in;
 reg local_bb2_cmp226_i217_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp296_i249_valid_out;
wire local_bb2_cmp296_i249_stall_in;
 reg local_bb2_cmp296_i249_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i250_valid_out;
wire local_bb2_cmp299_i250_stall_in;
 reg local_bb2_cmp299_i250_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i250_inputs_ready;
wire local_bb2_cmp299_i250_stall_local;
wire local_bb2_cmp299_i250;

assign local_bb2_cmp299_i250_inputs_ready = (rnode_173to175_bb2_shr16_i93_0_valid_out_NO_SHIFT_REG & rnode_173to175_bb2_cmp37_i105_0_valid_out_2_NO_SHIFT_REG & rnode_173to175_bb2_and17_i94_0_valid_out_NO_SHIFT_REG & rnode_173to175_bb2_cmp37_i105_0_valid_out_0_NO_SHIFT_REG & rnode_174to175_bb2_and193_i183_0_valid_out_2_NO_SHIFT_REG & rnode_173to175_bb2_cmp37_i105_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2_and195_i184_0_valid_out_NO_SHIFT_REG & rnode_174to175_bb2_and193_i183_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2_and198_i185_0_valid_out_NO_SHIFT_REG & rnode_174to175_bb2_and193_i183_0_valid_out_0_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i198_0_valid_out_1_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i198_0_valid_out_2_NO_SHIFT_REG & rnode_174to175_bb2__and_i_i198_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_cmp299_i250 = (local_bb2_and270_i234 == 32'h4);
assign local_bb2_and269_i237_valid_out = 1'b1;
assign local_bb2_add245_i223_valid_out = 1'b1;
assign local_bb2_notrhs_i228_valid_out = 1'b1;
assign local_bb2_not_cmp37_i211_valid_out_1 = 1'b1;
assign local_bb2_shr271_i235_valid_out = 1'b1;
assign local_bb2_cmp226_i217_valid_out = 1'b1;
assign local_bb2_cmp296_i249_valid_out = 1'b1;
assign local_bb2_cmp299_i250_valid_out = 1'b1;
assign rnode_173to175_bb2_shr16_i93_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp37_i105_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_and17_i94_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp37_i105_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and193_i183_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_173to175_bb2_cmp37_i105_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and195_i184_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and193_i183_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and198_i185_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2_and193_i183_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i198_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i198_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_174to175_bb2__and_i_i198_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_and269_i237_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add245_i223_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_notrhs_i228_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_not_cmp37_i211_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr271_i235_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp226_i217_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp296_i249_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp299_i250_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_and269_i237_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i250_inputs_ready & (local_bb2_and269_i237_consumed_0_NO_SHIFT_REG | ~(local_bb2_and269_i237_stall_in)) & local_bb2_cmp299_i250_stall_local);
		local_bb2_add245_i223_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i250_inputs_ready & (local_bb2_add245_i223_consumed_0_NO_SHIFT_REG | ~(local_bb2_add245_i223_stall_in)) & local_bb2_cmp299_i250_stall_local);
		local_bb2_notrhs_i228_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i250_inputs_ready & (local_bb2_notrhs_i228_consumed_0_NO_SHIFT_REG | ~(local_bb2_notrhs_i228_stall_in)) & local_bb2_cmp299_i250_stall_local);
		local_bb2_not_cmp37_i211_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp299_i250_inputs_ready & (local_bb2_not_cmp37_i211_consumed_1_NO_SHIFT_REG | ~(local_bb2_not_cmp37_i211_stall_in_1)) & local_bb2_cmp299_i250_stall_local);
		local_bb2_shr271_i235_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i250_inputs_ready & (local_bb2_shr271_i235_consumed_0_NO_SHIFT_REG | ~(local_bb2_shr271_i235_stall_in)) & local_bb2_cmp299_i250_stall_local);
		local_bb2_cmp226_i217_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i250_inputs_ready & (local_bb2_cmp226_i217_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp226_i217_stall_in)) & local_bb2_cmp299_i250_stall_local);
		local_bb2_cmp296_i249_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i250_inputs_ready & (local_bb2_cmp296_i249_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp296_i249_stall_in)) & local_bb2_cmp299_i250_stall_local);
		local_bb2_cmp299_i250_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i250_inputs_ready & (local_bb2_cmp299_i250_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp299_i250_stall_in)) & local_bb2_cmp299_i250_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_and270_i718_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i718_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and270_i718_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i718_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and270_i718_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i718_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i718_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and270_i718_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_and270_i718_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_and270_i718_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_and270_i718_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_and270_i718_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_and270_i718_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_and270_i718),
	.data_out(rnode_175to176_bb2_and270_i718_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_and270_i718_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_and270_i718_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_and270_i718_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_and270_i718_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_and270_i718_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and270_i718_stall_in = 1'b0;
assign rnode_175to176_bb2_and270_i718_0_NO_SHIFT_REG = rnode_175to176_bb2_and270_i718_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_and270_i718_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and270_i718_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_add246_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add246_i_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add246_i_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add246_i_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_add246_i_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_add246_i_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_add246_i_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_add246_i_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_add246_i_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_add246_i),
	.data_out(rnode_175to176_bb2_add246_i_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_add246_i_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_add246_i_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_add246_i_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_add246_i_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_add246_i_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add246_i_stall_in_1 = 1'b0;
assign rnode_175to176_bb2_add246_i_0_NO_SHIFT_REG = rnode_175to176_bb2_add246_i_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_add246_i_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add246_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_not__46_i716_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not__46_i716_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not__46_i716_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not__46_i716_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not__46_i716_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not__46_i716_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not__46_i716_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not__46_i716_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_not__46_i716_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_not__46_i716_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_not__46_i716_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_not__46_i716_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_not__46_i716_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_not__46_i716),
	.data_out(rnode_175to176_bb2_not__46_i716_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_not__46_i716_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_not__46_i716_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_not__46_i716_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_not__46_i716_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_not__46_i716_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not__46_i716_stall_in = 1'b0;
assign rnode_175to176_bb2_not__46_i716_0_NO_SHIFT_REG = rnode_175to176_bb2_not__46_i716_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_not__46_i716_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not__46_i716_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_not_cmp38_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp38_i_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_not_cmp38_i_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_not_cmp38_i_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_not_cmp38_i_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_not_cmp38_i_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_not_cmp38_i_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_not_cmp38_i),
	.data_out(rnode_175to176_bb2_not_cmp38_i_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_not_cmp38_i_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_not_cmp38_i_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_not_cmp38_i_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_not_cmp38_i_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_not_cmp38_i_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not_cmp38_i_stall_in_1 = 1'b0;
assign rnode_175to176_bb2_not_cmp38_i_0_NO_SHIFT_REG = rnode_175to176_bb2_not_cmp38_i_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_not_cmp38_i_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not_cmp38_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_shr272_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_shr272_i_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_shr272_i_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr272_i_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_shr272_i_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_shr272_i_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_shr272_i_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_shr272_i_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_shr272_i_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_shr272_i),
	.data_out(rnode_175to176_bb2_shr272_i_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_shr272_i_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_shr272_i_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_shr272_i_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_shr272_i_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_shr272_i_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr272_i_stall_in = 1'b0;
assign rnode_175to176_bb2_shr272_i_0_NO_SHIFT_REG = rnode_175to176_bb2_shr272_i_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_shr272_i_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_shr272_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp227_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp227_i_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp227_i_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp227_i_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp227_i_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp227_i_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp227_i_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp227_i),
	.data_out(rnode_175to176_bb2_cmp227_i_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp227_i_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp227_i_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp227_i_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp227_i_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp227_i_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp227_i_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp227_i_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp227_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_cmp227_i_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp227_i_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp227_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_cmp227_i_1_NO_SHIFT_REG = rnode_175to176_bb2_cmp227_i_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp297_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp297_i_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp297_i_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp297_i_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp297_i_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp297_i_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp297_i_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp297_i),
	.data_out(rnode_175to176_bb2_cmp297_i_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp297_i_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp297_i_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp297_i_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp297_i_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp297_i_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp297_i_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp297_i_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp297_i_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp297_i_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp297_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp300_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp300_i_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp300_i_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp300_i_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp300_i_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp300_i_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp300_i_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp300_i),
	.data_out(rnode_175to176_bb2_cmp300_i_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp300_i_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp300_i_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp300_i_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp300_i_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp300_i_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp300_i_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp300_i_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp300_i_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp300_i_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp300_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shl274_i1799_stall_local;
wire [31:0] local_bb2_shl274_i1799;

assign local_bb2_shl274_i1799 = (rnode_175to176_bb2_and270_i1798_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and248_i1785_stall_local;
wire [31:0] local_bb2_and248_i1785;

assign local_bb2_and248_i1785 = (rnode_175to176_bb2_add246_i1784_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp259_i1792_stall_local;
wire local_bb2_cmp259_i1792;

assign local_bb2_cmp259_i1792 = ($signed(rnode_175to176_bb2_add246_i1784_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb2_and273_i1797_stall_local;
wire [31:0] local_bb2_and273_i1797;

assign local_bb2_and273_i1797 = (rnode_175to176_bb2_shr272_i1796_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp227_not_i1779_stall_local;
wire local_bb2_cmp227_not_i1779;

assign local_bb2_cmp227_not_i1779 = (rnode_175to176_bb2_cmp227_i1778_0_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp29749_i1814_stall_local;
wire [31:0] local_bb2_cmp29749_i1814;

assign local_bb2_cmp29749_i1814[31:1] = 31'h0;
assign local_bb2_cmp29749_i1814[0] = rnode_175to176_bb2_cmp297_i1810_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_conv301_i1812_stall_local;
wire [31:0] local_bb2_conv301_i1812;

assign local_bb2_conv301_i1812[31:1] = 31'h0;
assign local_bb2_conv301_i1812[0] = rnode_175to176_bb2_cmp300_i1811_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_and269_i1249_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i1249_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and269_i1249_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i1249_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and269_i1249_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i1249_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i1249_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i1249_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_and269_i1249_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_and269_i1249_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_and269_i1249_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_and269_i1249_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_and269_i1249_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_and269_i1249),
	.data_out(rnode_175to176_bb2_and269_i1249_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_and269_i1249_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_and269_i1249_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_and269_i1249_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_and269_i1249_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_and269_i1249_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and269_i1249_stall_in = 1'b0;
assign rnode_175to176_bb2_and269_i1249_0_NO_SHIFT_REG = rnode_175to176_bb2_and269_i1249_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_and269_i1249_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and269_i1249_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_add245_i1235_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i1235_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add245_i1235_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i1235_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i1235_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add245_i1235_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i1235_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add245_i1235_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i1235_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i1235_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i1235_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_add245_i1235_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_add245_i1235_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_add245_i1235_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_add245_i1235_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_add245_i1235_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_add245_i1235),
	.data_out(rnode_175to176_bb2_add245_i1235_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_add245_i1235_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_add245_i1235_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_add245_i1235_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_add245_i1235_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_add245_i1235_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add245_i1235_stall_in = 1'b0;
assign rnode_175to176_bb2_add245_i1235_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add245_i1235_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_add245_i1235_0_NO_SHIFT_REG = rnode_175to176_bb2_add245_i1235_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_add245_i1235_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_add245_i1235_1_NO_SHIFT_REG = rnode_175to176_bb2_add245_i1235_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_notrhs_i1240_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1240_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1240_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1240_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1240_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1240_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1240_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i1240_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_notrhs_i1240_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_notrhs_i1240_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_notrhs_i1240_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_notrhs_i1240_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_notrhs_i1240_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_notrhs_i1240),
	.data_out(rnode_175to176_bb2_notrhs_i1240_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_notrhs_i1240_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_notrhs_i1240_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_notrhs_i1240_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_notrhs_i1240_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_notrhs_i1240_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_notrhs_i1240_stall_in = 1'b0;
assign rnode_175to176_bb2_notrhs_i1240_0_NO_SHIFT_REG = rnode_175to176_bb2_notrhs_i1240_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_notrhs_i1240_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_notrhs_i1240_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_not_cmp37_i1223_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i1223_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i1223_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i1223_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i1223_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i1223_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_not_cmp37_i1223_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_not_cmp37_i1223_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_not_cmp37_i1223_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_not_cmp37_i1223),
	.data_out(rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not_cmp37_i1223_stall_in_1 = 1'b0;
assign rnode_175to176_bb2_not_cmp37_i1223_0_NO_SHIFT_REG = rnode_175to176_bb2_not_cmp37_i1223_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_not_cmp37_i1223_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not_cmp37_i1223_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_shr271_i1247_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i1247_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_shr271_i1247_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i1247_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_shr271_i1247_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i1247_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i1247_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i1247_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_shr271_i1247_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_shr271_i1247_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_shr271_i1247_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_shr271_i1247_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_shr271_i1247_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_shr271_i1247),
	.data_out(rnode_175to176_bb2_shr271_i1247_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_shr271_i1247_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_shr271_i1247_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_shr271_i1247_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_shr271_i1247_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_shr271_i1247_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr271_i1247_stall_in = 1'b0;
assign rnode_175to176_bb2_shr271_i1247_0_NO_SHIFT_REG = rnode_175to176_bb2_shr271_i1247_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_shr271_i1247_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_shr271_i1247_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp226_i1229_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i1229_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp226_i1229_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp226_i1229_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp226_i1229_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp226_i1229_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp226_i1229_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp226_i1229),
	.data_out(rnode_175to176_bb2_cmp226_i1229_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp226_i1229_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp226_i1229_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp226_i1229_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp226_i1229_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp226_i1229_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp226_i1229_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp226_i1229_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp226_i1229_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_cmp226_i1229_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp226_i1229_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp226_i1229_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_cmp226_i1229_1_NO_SHIFT_REG = rnode_175to176_bb2_cmp226_i1229_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp296_i1261_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i1261_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i1261_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i1261_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i1261_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i1261_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i1261_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i1261_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp296_i1261_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp296_i1261_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp296_i1261_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp296_i1261_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp296_i1261_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp296_i1261),
	.data_out(rnode_175to176_bb2_cmp296_i1261_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp296_i1261_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp296_i1261_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp296_i1261_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp296_i1261_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp296_i1261_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp296_i1261_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp296_i1261_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp296_i1261_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp296_i1261_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp296_i1261_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp299_i1262_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i1262_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i1262_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i1262_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i1262_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i1262_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i1262_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i1262_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp299_i1262_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp299_i1262_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp299_i1262_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp299_i1262_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp299_i1262_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp299_i1262),
	.data_out(rnode_175to176_bb2_cmp299_i1262_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp299_i1262_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp299_i1262_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp299_i1262_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp299_i1262_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp299_i1262_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp299_i1262_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp299_i1262_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp299_i1262_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp299_i1262_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp299_i1262_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_and269_i237_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i237_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and269_i237_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i237_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_and269_i237_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i237_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i237_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_and269_i237_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_and269_i237_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_and269_i237_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_and269_i237_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_and269_i237_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_and269_i237_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_and269_i237),
	.data_out(rnode_175to176_bb2_and269_i237_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_and269_i237_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_and269_i237_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_and269_i237_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_and269_i237_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_and269_i237_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and269_i237_stall_in = 1'b0;
assign rnode_175to176_bb2_and269_i237_0_NO_SHIFT_REG = rnode_175to176_bb2_and269_i237_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_and269_i237_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and269_i237_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_add245_i223_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i223_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add245_i223_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i223_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i223_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add245_i223_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i223_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_add245_i223_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i223_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i223_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_add245_i223_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_add245_i223_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_add245_i223_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_add245_i223_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_add245_i223_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_add245_i223_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_add245_i223),
	.data_out(rnode_175to176_bb2_add245_i223_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_add245_i223_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_add245_i223_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_add245_i223_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_add245_i223_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_add245_i223_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add245_i223_stall_in = 1'b0;
assign rnode_175to176_bb2_add245_i223_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add245_i223_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_add245_i223_0_NO_SHIFT_REG = rnode_175to176_bb2_add245_i223_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_add245_i223_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_add245_i223_1_NO_SHIFT_REG = rnode_175to176_bb2_add245_i223_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_notrhs_i228_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i228_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i228_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i228_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i228_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i228_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i228_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_notrhs_i228_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_notrhs_i228_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_notrhs_i228_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_notrhs_i228_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_notrhs_i228_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_notrhs_i228_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_notrhs_i228),
	.data_out(rnode_175to176_bb2_notrhs_i228_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_notrhs_i228_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_notrhs_i228_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_notrhs_i228_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_notrhs_i228_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_notrhs_i228_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_notrhs_i228_stall_in = 1'b0;
assign rnode_175to176_bb2_notrhs_i228_0_NO_SHIFT_REG = rnode_175to176_bb2_notrhs_i228_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_notrhs_i228_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_notrhs_i228_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_not_cmp37_i211_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i211_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i211_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i211_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i211_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i211_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i211_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_not_cmp37_i211_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_not_cmp37_i211_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_not_cmp37_i211_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_not_cmp37_i211_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_not_cmp37_i211_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_not_cmp37_i211_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_not_cmp37_i211),
	.data_out(rnode_175to176_bb2_not_cmp37_i211_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_not_cmp37_i211_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_not_cmp37_i211_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_not_cmp37_i211_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_not_cmp37_i211_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_not_cmp37_i211_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not_cmp37_i211_stall_in_1 = 1'b0;
assign rnode_175to176_bb2_not_cmp37_i211_0_NO_SHIFT_REG = rnode_175to176_bb2_not_cmp37_i211_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_not_cmp37_i211_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not_cmp37_i211_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_shr271_i235_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i235_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_shr271_i235_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i235_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_175to176_bb2_shr271_i235_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i235_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i235_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_shr271_i235_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_shr271_i235_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_shr271_i235_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_shr271_i235_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_shr271_i235_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_shr271_i235_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_shr271_i235),
	.data_out(rnode_175to176_bb2_shr271_i235_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_shr271_i235_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_shr271_i235_0_reg_176_fifo.DATA_WIDTH = 32;
defparam rnode_175to176_bb2_shr271_i235_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_shr271_i235_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_shr271_i235_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr271_i235_stall_in = 1'b0;
assign rnode_175to176_bb2_shr271_i235_0_NO_SHIFT_REG = rnode_175to176_bb2_shr271_i235_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_shr271_i235_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_shr271_i235_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp226_i217_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_1_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_valid_out_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_stall_in_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp226_i217_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp226_i217_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp226_i217_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp226_i217_0_stall_in_0_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp226_i217_0_valid_out_0_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp226_i217_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp226_i217),
	.data_out(rnode_175to176_bb2_cmp226_i217_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp226_i217_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp226_i217_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp226_i217_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp226_i217_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp226_i217_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp226_i217_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp226_i217_0_stall_in_0_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp226_i217_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_cmp226_i217_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp226_i217_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp226_i217_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_175to176_bb2_cmp226_i217_1_NO_SHIFT_REG = rnode_175to176_bb2_cmp226_i217_0_reg_176_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp296_i249_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i249_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i249_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i249_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i249_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i249_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i249_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp296_i249_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp296_i249_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp296_i249_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp296_i249_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp296_i249_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp296_i249_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp296_i249),
	.data_out(rnode_175to176_bb2_cmp296_i249_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp296_i249_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp296_i249_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp296_i249_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp296_i249_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp296_i249_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp296_i249_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp296_i249_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp296_i249_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp296_i249_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp296_i249_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_175to176_bb2_cmp299_i250_0_valid_out_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i250_0_stall_in_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i250_0_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i250_0_reg_176_inputs_ready_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i250_0_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i250_0_valid_out_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i250_0_stall_in_reg_176_NO_SHIFT_REG;
 logic rnode_175to176_bb2_cmp299_i250_0_stall_out_reg_176_NO_SHIFT_REG;

acl_data_fifo rnode_175to176_bb2_cmp299_i250_0_reg_176_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_175to176_bb2_cmp299_i250_0_reg_176_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_175to176_bb2_cmp299_i250_0_stall_in_reg_176_NO_SHIFT_REG),
	.valid_out(rnode_175to176_bb2_cmp299_i250_0_valid_out_reg_176_NO_SHIFT_REG),
	.stall_out(rnode_175to176_bb2_cmp299_i250_0_stall_out_reg_176_NO_SHIFT_REG),
	.data_in(local_bb2_cmp299_i250),
	.data_out(rnode_175to176_bb2_cmp299_i250_0_reg_176_NO_SHIFT_REG)
);

defparam rnode_175to176_bb2_cmp299_i250_0_reg_176_fifo.DEPTH = 1;
defparam rnode_175to176_bb2_cmp299_i250_0_reg_176_fifo.DATA_WIDTH = 1;
defparam rnode_175to176_bb2_cmp299_i250_0_reg_176_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_175to176_bb2_cmp299_i250_0_reg_176_fifo.IMPL = "shift_reg";

assign rnode_175to176_bb2_cmp299_i250_0_reg_176_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp299_i250_stall_in = 1'b0;
assign rnode_175to176_bb2_cmp299_i250_0_NO_SHIFT_REG = rnode_175to176_bb2_cmp299_i250_0_reg_176_NO_SHIFT_REG;
assign rnode_175to176_bb2_cmp299_i250_0_stall_in_reg_176_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp299_i250_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shl274_i_stall_local;
wire [31:0] local_bb2_shl274_i;

assign local_bb2_shl274_i = (rnode_175to176_bb2_and270_i718_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp259_i_stall_local;
wire local_bb2_cmp259_i;

assign local_bb2_cmp259_i = ($signed(rnode_175to176_bb2_add246_i_0_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb2_and273_i_stall_local;
wire [31:0] local_bb2_and273_i;

assign local_bb2_and273_i = (rnode_175to176_bb2_shr272_i_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp227_not_i_stall_local;
wire local_bb2_cmp227_not_i;

assign local_bb2_cmp227_not_i = (rnode_175to176_bb2_cmp227_i_0_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__47_i717_stall_local;
wire local_bb2__47_i717;

assign local_bb2__47_i717 = (rnode_175to176_bb2_cmp227_i_1_NO_SHIFT_REG | rnode_175to176_bb2_not__46_i716_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp29749_i_stall_local;
wire [31:0] local_bb2_cmp29749_i;

assign local_bb2_cmp29749_i[31:1] = 31'h0;
assign local_bb2_cmp29749_i[0] = rnode_175to176_bb2_cmp297_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_conv301_i_stall_local;
wire [31:0] local_bb2_conv301_i;

assign local_bb2_conv301_i[31:1] = 31'h0;
assign local_bb2_conv301_i[0] = rnode_175to176_bb2_cmp300_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_notlhs_i1788_stall_local;
wire local_bb2_notlhs_i1788;

assign local_bb2_notlhs_i1788 = (local_bb2_and248_i1785 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or275_i1800_stall_local;
wire [31:0] local_bb2_or275_i1800;

assign local_bb2_or275_i1800 = (local_bb2_and273_i1797 | local_bb2_shl274_i1799);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge12_i1780_stall_local;
wire local_bb2_brmerge12_i1780;

assign local_bb2_brmerge12_i1780 = (local_bb2_cmp227_not_i1779 | rnode_175to176_bb2_not_cmp38_i1772_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot263__i1793_stall_local;
wire local_bb2_lnot263__i1793;

assign local_bb2_lnot263__i1793 = (local_bb2_cmp259_i1792 & local_bb2_cmp227_not_i1779);

// This section implements an unregistered operation.
// 
wire local_bb2_shl273_i1250_stall_local;
wire [31:0] local_bb2_shl273_i1250;

assign local_bb2_shl273_i1250 = (rnode_175to176_bb2_and269_i1249_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and247_i1236_stall_local;
wire [31:0] local_bb2_and247_i1236;

assign local_bb2_and247_i1236 = (rnode_175to176_bb2_add245_i1235_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp258_i1243_stall_local;
wire local_bb2_cmp258_i1243;

assign local_bb2_cmp258_i1243 = ($signed(rnode_175to176_bb2_add245_i1235_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb2_and272_i1248_stall_local;
wire [31:0] local_bb2_and272_i1248;

assign local_bb2_and272_i1248 = (rnode_175to176_bb2_shr271_i1247_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_not_i1230_stall_local;
wire local_bb2_cmp226_not_i1230;

assign local_bb2_cmp226_not_i1230 = (rnode_175to176_bb2_cmp226_i1229_0_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp29649_i1265_stall_local;
wire [31:0] local_bb2_cmp29649_i1265;

assign local_bb2_cmp29649_i1265[31:1] = 31'h0;
assign local_bb2_cmp29649_i1265[0] = rnode_175to176_bb2_cmp296_i1261_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_conv300_i1263_stall_local;
wire [31:0] local_bb2_conv300_i1263;

assign local_bb2_conv300_i1263[31:1] = 31'h0;
assign local_bb2_conv300_i1263[0] = rnode_175to176_bb2_cmp299_i1262_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shl273_i238_stall_local;
wire [31:0] local_bb2_shl273_i238;

assign local_bb2_shl273_i238 = (rnode_175to176_bb2_and269_i237_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_and247_i224_stall_local;
wire [31:0] local_bb2_and247_i224;

assign local_bb2_and247_i224 = (rnode_175to176_bb2_add245_i223_0_NO_SHIFT_REG & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp258_i231_stall_local;
wire local_bb2_cmp258_i231;

assign local_bb2_cmp258_i231 = ($signed(rnode_175to176_bb2_add245_i223_1_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb2_and272_i236_stall_local;
wire [31:0] local_bb2_and272_i236;

assign local_bb2_and272_i236 = (rnode_175to176_bb2_shr271_i235_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_not_i218_stall_local;
wire local_bb2_cmp226_not_i218;

assign local_bb2_cmp226_not_i218 = (rnode_175to176_bb2_cmp226_i217_0_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp29649_i253_stall_local;
wire [31:0] local_bb2_cmp29649_i253;

assign local_bb2_cmp29649_i253[31:1] = 31'h0;
assign local_bb2_cmp29649_i253[0] = rnode_175to176_bb2_cmp296_i249_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_conv300_i251_stall_local;
wire [31:0] local_bb2_conv300_i251;

assign local_bb2_conv300_i251[31:1] = 31'h0;
assign local_bb2_conv300_i251[0] = rnode_175to176_bb2_cmp299_i250_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_or275_i719_stall_local;
wire [31:0] local_bb2_or275_i719;

assign local_bb2_or275_i719 = (local_bb2_and273_i | local_bb2_shl274_i);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge12_i711_stall_local;
wire local_bb2_brmerge12_i711;

assign local_bb2_brmerge12_i711 = (local_bb2_cmp227_not_i | rnode_175to176_bb2_not_cmp38_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot263__i_stall_local;
wire local_bb2_lnot263__i;

assign local_bb2_lnot263__i = (local_bb2_cmp259_i & local_bb2_cmp227_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u128_stall_local;
wire [31:0] local_bb2_var__u128;

assign local_bb2_var__u128[31:1] = 31'h0;
assign local_bb2_var__u128[0] = local_bb2__47_i717;

// This section implements an unregistered operation.
// 
wire local_bb2_not__46_i1790_stall_local;
wire local_bb2_not__46_i1790;

assign local_bb2_not__46_i1790 = (rnode_175to176_bb2_notrhs_i1789_0_NO_SHIFT_REG | local_bb2_notlhs_i1788);

// This section implements an unregistered operation.
// 
wire local_bb2_resultSign_0_i1781_stall_local;
wire [31:0] local_bb2_resultSign_0_i1781;

assign local_bb2_resultSign_0_i1781 = (local_bb2_brmerge12_i1780 ? rnode_175to176_bb2_and35_i1664_0_NO_SHIFT_REG : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or2672_i1794_stall_local;
wire local_bb2_or2672_i1794;

assign local_bb2_or2672_i1794 = (rnode_175to176_bb2_var__u102_0_NO_SHIFT_REG | local_bb2_lnot263__i1793);

// This section implements an unregistered operation.
// 
wire local_bb2_notlhs_i1239_stall_local;
wire local_bb2_notlhs_i1239;

assign local_bb2_notlhs_i1239 = (local_bb2_and247_i1236 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or274_i1251_stall_local;
wire [31:0] local_bb2_or274_i1251;

assign local_bb2_or274_i1251 = (local_bb2_and272_i1248 | local_bb2_shl273_i1250);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge12_i1231_stall_local;
wire local_bb2_brmerge12_i1231;

assign local_bb2_brmerge12_i1231 = (local_bb2_cmp226_not_i1230 | rnode_175to176_bb2_not_cmp37_i1223_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot262__i1244_stall_local;
wire local_bb2_lnot262__i1244;

assign local_bb2_lnot262__i1244 = (local_bb2_cmp258_i1243 & local_bb2_cmp226_not_i1230);

// This section implements an unregistered operation.
// 
wire local_bb2_notlhs_i227_stall_local;
wire local_bb2_notlhs_i227;

assign local_bb2_notlhs_i227 = (local_bb2_and247_i224 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or274_i239_stall_local;
wire [31:0] local_bb2_or274_i239;

assign local_bb2_or274_i239 = (local_bb2_and272_i236 | local_bb2_shl273_i238);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge12_i219_stall_local;
wire local_bb2_brmerge12_i219;

assign local_bb2_brmerge12_i219 = (local_bb2_cmp226_not_i218 | rnode_175to176_bb2_not_cmp37_i211_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot262__i232_stall_local;
wire local_bb2_lnot262__i232;

assign local_bb2_lnot262__i232 = (local_bb2_cmp258_i231 & local_bb2_cmp226_not_i218);

// This section implements an unregistered operation.
// 
wire local_bb2_resultSign_0_i712_stall_local;
wire [31:0] local_bb2_resultSign_0_i712;

assign local_bb2_resultSign_0_i712 = (local_bb2_brmerge12_i711 ? rnode_175to176_bb2_and35_i652_0_NO_SHIFT_REG : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or2672_i_stall_local;
wire local_bb2_or2672_i;

assign local_bb2_or2672_i = (rnode_175to176_bb2_var__u107_0_NO_SHIFT_REG | local_bb2_lnot263__i);

// This section implements an unregistered operation.
// 
wire local_bb2__47_i1791_stall_local;
wire local_bb2__47_i1791;

assign local_bb2__47_i1791 = (rnode_175to176_bb2_cmp227_i1778_1_NO_SHIFT_REG | local_bb2_not__46_i1790);

// This section implements an unregistered operation.
// 
wire local_bb2_or276_i1801_stall_local;
wire [31:0] local_bb2_or276_i1801;

assign local_bb2_or276_i1801 = (local_bb2_or275_i1800 | local_bb2_resultSign_0_i1781);

// This section implements an unregistered operation.
// 
wire local_bb2_or2885_i1804_stall_local;
wire local_bb2_or2885_i1804;

assign local_bb2_or2885_i1804 = (local_bb2_or2672_i1794 | rnode_175to176_bb2__26_i1679_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u129_stall_local;
wire [31:0] local_bb2_var__u129;

assign local_bb2_var__u129[31:1] = 31'h0;
assign local_bb2_var__u129[0] = local_bb2_or2672_i1794;

// This section implements an unregistered operation.
// 
wire local_bb2_not__46_i1241_stall_local;
wire local_bb2_not__46_i1241;

assign local_bb2_not__46_i1241 = (rnode_175to176_bb2_notrhs_i1240_0_NO_SHIFT_REG | local_bb2_notlhs_i1239);

// This section implements an unregistered operation.
// 
wire local_bb2_resultSign_0_i1232_stall_local;
wire [31:0] local_bb2_resultSign_0_i1232;

assign local_bb2_resultSign_0_i1232 = (local_bb2_brmerge12_i1231 ? rnode_175to176_bb2_and35_i1115_0_NO_SHIFT_REG : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or2662_i1245_stall_local;
wire local_bb2_or2662_i1245;

assign local_bb2_or2662_i1245 = (rnode_175to176_bb2_var__u111_0_NO_SHIFT_REG | local_bb2_lnot262__i1244);

// This section implements an unregistered operation.
// 
wire local_bb2_not__46_i229_stall_local;
wire local_bb2_not__46_i229;

assign local_bb2_not__46_i229 = (rnode_175to176_bb2_notrhs_i228_0_NO_SHIFT_REG | local_bb2_notlhs_i227);

// This section implements an unregistered operation.
// 
wire local_bb2_resultSign_0_i220_stall_local;
wire [31:0] local_bb2_resultSign_0_i220;

assign local_bb2_resultSign_0_i220 = (local_bb2_brmerge12_i219 ? rnode_175to176_bb2_and35_i103_0_NO_SHIFT_REG : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or2662_i233_stall_local;
wire local_bb2_or2662_i233;

assign local_bb2_or2662_i233 = (rnode_175to176_bb2_var__u114_0_NO_SHIFT_REG | local_bb2_lnot262__i232);

// This section implements an unregistered operation.
// 
wire local_bb2_or276_i_stall_local;
wire [31:0] local_bb2_or276_i;

assign local_bb2_or276_i = (local_bb2_or275_i719 | local_bb2_resultSign_0_i712);

// This section implements an unregistered operation.
// 
wire local_bb2_or2814_i_stall_local;
wire local_bb2_or2814_i;

assign local_bb2_or2814_i = (local_bb2__47_i717 | local_bb2_or2672_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or2885_i_stall_local;
wire local_bb2_or2885_i;

assign local_bb2_or2885_i = (local_bb2_or2672_i | rnode_175to176_bb2__26_i665_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u130_stall_local;
wire [31:0] local_bb2_var__u130;

assign local_bb2_var__u130[31:1] = 31'h0;
assign local_bb2_var__u130[0] = local_bb2_or2672_i;

// This section implements an unregistered operation.
// 
wire local_bb2_or2814_i1802_stall_local;
wire local_bb2_or2814_i1802;

assign local_bb2_or2814_i1802 = (local_bb2__47_i1791 | local_bb2_or2672_i1794);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u131_stall_local;
wire [31:0] local_bb2_var__u131;

assign local_bb2_var__u131[31:1] = 31'h0;
assign local_bb2_var__u131[0] = local_bb2__47_i1791;

// This section implements an unregistered operation.
// 
wire local_bb2_cond290_i1805_stall_local;
wire [31:0] local_bb2_cond290_i1805;

assign local_bb2_cond290_i1805 = (local_bb2_or2885_i1804 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext311_i1817_stall_local;
wire [31:0] local_bb2_lnot_ext311_i1817;

assign local_bb2_lnot_ext311_i1817 = (local_bb2_var__u129 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__47_i1242_stall_local;
wire local_bb2__47_i1242;

assign local_bb2__47_i1242 = (rnode_175to176_bb2_cmp226_i1229_1_NO_SHIFT_REG | local_bb2_not__46_i1241);

// This section implements an unregistered operation.
// 
wire local_bb2_or275_i1252_stall_local;
wire [31:0] local_bb2_or275_i1252;

assign local_bb2_or275_i1252 = (local_bb2_or274_i1251 | local_bb2_resultSign_0_i1232);

// This section implements an unregistered operation.
// 
wire local_bb2_or2875_i1255_stall_local;
wire local_bb2_or2875_i1255;

assign local_bb2_or2875_i1255 = (local_bb2_or2662_i1245 | rnode_175to176_bb2__26_i1130_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u132_stall_local;
wire [31:0] local_bb2_var__u132;

assign local_bb2_var__u132[31:1] = 31'h0;
assign local_bb2_var__u132[0] = local_bb2_or2662_i1245;

// This section implements an unregistered operation.
// 
wire local_bb2__47_i230_stall_local;
wire local_bb2__47_i230;

assign local_bb2__47_i230 = (rnode_175to176_bb2_cmp226_i217_1_NO_SHIFT_REG | local_bb2_not__46_i229);

// This section implements an unregistered operation.
// 
wire local_bb2_or275_i240_stall_local;
wire [31:0] local_bb2_or275_i240;

assign local_bb2_or275_i240 = (local_bb2_or274_i239 | local_bb2_resultSign_0_i220);

// This section implements an unregistered operation.
// 
wire local_bb2_or2875_i243_stall_local;
wire local_bb2_or2875_i243;

assign local_bb2_or2875_i243 = (local_bb2_or2662_i233 | rnode_175to176_bb2__26_i118_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u133_stall_local;
wire [31:0] local_bb2_var__u133;

assign local_bb2_var__u133[31:1] = 31'h0;
assign local_bb2_var__u133[0] = local_bb2_or2662_i233;

// This section implements an unregistered operation.
// 
wire local_bb2_cond283_i_stall_local;
wire [31:0] local_bb2_cond283_i;

assign local_bb2_cond283_i = (local_bb2_or2814_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond290_i_stall_local;
wire [31:0] local_bb2_cond290_i;

assign local_bb2_cond290_i = (local_bb2_or2885_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext311_i_stall_local;
wire [31:0] local_bb2_lnot_ext311_i;

assign local_bb2_lnot_ext311_i = (local_bb2_var__u130 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cond283_i1803_stall_local;
wire [31:0] local_bb2_cond283_i1803;

assign local_bb2_cond283_i1803 = (local_bb2_or2814_i1802 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i1808_stall_local;
wire [31:0] local_bb2_or295_i1808;

assign local_bb2_or295_i1808 = (local_bb2_cond290_i1805 | local_bb2_cond293_i1806);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i1819_stall_local;
wire [31:0] local_bb2_reduction_0_i1819;

assign local_bb2_reduction_0_i1819 = (local_bb2_lnot_ext311_i1817 & local_bb2_lnot_ext_i1816);

// This section implements an unregistered operation.
// 
wire local_bb2_or2804_i1253_stall_local;
wire local_bb2_or2804_i1253;

assign local_bb2_or2804_i1253 = (local_bb2__47_i1242 | local_bb2_or2662_i1245);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u134_stall_local;
wire [31:0] local_bb2_var__u134;

assign local_bb2_var__u134[31:1] = 31'h0;
assign local_bb2_var__u134[0] = local_bb2__47_i1242;

// This section implements an unregistered operation.
// 
wire local_bb2_cond289_i1256_stall_local;
wire [31:0] local_bb2_cond289_i1256;

assign local_bb2_cond289_i1256 = (local_bb2_or2875_i1255 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext310_i1268_stall_local;
wire [31:0] local_bb2_lnot_ext310_i1268;

assign local_bb2_lnot_ext310_i1268 = (local_bb2_var__u132 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or2804_i241_stall_local;
wire local_bb2_or2804_i241;

assign local_bb2_or2804_i241 = (local_bb2__47_i230 | local_bb2_or2662_i233);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u135_stall_local;
wire [31:0] local_bb2_var__u135;

assign local_bb2_var__u135[31:1] = 31'h0;
assign local_bb2_var__u135[0] = local_bb2__47_i230;

// This section implements an unregistered operation.
// 
wire local_bb2_cond289_i244_stall_local;
wire [31:0] local_bb2_cond289_i244;

assign local_bb2_cond289_i244 = (local_bb2_or2875_i243 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext310_i256_stall_local;
wire [31:0] local_bb2_lnot_ext310_i256;

assign local_bb2_lnot_ext310_i256 = (local_bb2_var__u133 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and294_i_stall_local;
wire [31:0] local_bb2_and294_i;

assign local_bb2_and294_i = (local_bb2_cond283_i & local_bb2_or276_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i720_stall_local;
wire [31:0] local_bb2_or295_i720;

assign local_bb2_or295_i720 = (local_bb2_cond290_i | local_bb2_cond293_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i723_stall_local;
wire [31:0] local_bb2_reduction_0_i723;

assign local_bb2_reduction_0_i723 = (local_bb2_lnot_ext311_i & local_bb2_lnot_ext_i722);

// This section implements an unregistered operation.
// 
wire local_bb2_and294_i1807_stall_local;
wire [31:0] local_bb2_and294_i1807;

assign local_bb2_and294_i1807 = (local_bb2_cond283_i1803 & local_bb2_or276_i1801);

// This section implements an unregistered operation.
// 
wire local_bb2_cond282_i1254_stall_local;
wire [31:0] local_bb2_cond282_i1254;

assign local_bb2_cond282_i1254 = (local_bb2_or2804_i1253 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or294_i1259_stall_local;
wire [31:0] local_bb2_or294_i1259;

assign local_bb2_or294_i1259 = (local_bb2_cond289_i1256 | local_bb2_cond292_i1257);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i1270_stall_local;
wire [31:0] local_bb2_reduction_0_i1270;

assign local_bb2_reduction_0_i1270 = (local_bb2_lnot_ext310_i1268 & local_bb2_lnot_ext_i1267);

// This section implements an unregistered operation.
// 
wire local_bb2_cond282_i242_stall_local;
wire [31:0] local_bb2_cond282_i242;

assign local_bb2_cond282_i242 = (local_bb2_or2804_i241 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or294_i247_stall_local;
wire [31:0] local_bb2_or294_i247;

assign local_bb2_or294_i247 = (local_bb2_cond289_i244 | local_bb2_cond292_i245);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i258_stall_local;
wire [31:0] local_bb2_reduction_0_i258;

assign local_bb2_reduction_0_i258 = (local_bb2_lnot_ext310_i256 & local_bb2_lnot_ext_i255);

// This section implements an unregistered operation.
// 
wire local_bb2_and303_i_stall_local;
wire [31:0] local_bb2_and303_i;

assign local_bb2_and303_i = (local_bb2_conv301_i & local_bb2_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or296_i_stall_local;
wire [31:0] local_bb2_or296_i;

assign local_bb2_or296_i = (local_bb2_or295_i720 | local_bb2_and294_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or296_i1809_stall_local;
wire [31:0] local_bb2_or296_i1809;

assign local_bb2_or296_i1809 = (local_bb2_or295_i1808 | local_bb2_and294_i1807);

// This section implements an unregistered operation.
// 
wire local_bb2_and303_i1813_stall_local;
wire [31:0] local_bb2_and303_i1813;

assign local_bb2_and303_i1813 = (local_bb2_conv301_i1812 & local_bb2_and294_i1807);

// This section implements an unregistered operation.
// 
wire local_bb2_and293_i1258_stall_local;
wire [31:0] local_bb2_and293_i1258;

assign local_bb2_and293_i1258 = (local_bb2_cond282_i1254 & local_bb2_or275_i1252);

// This section implements an unregistered operation.
// 
wire local_bb2_and293_i246_stall_local;
wire [31:0] local_bb2_and293_i246;

assign local_bb2_and293_i246 = (local_bb2_cond282_i242 & local_bb2_or275_i240);

// This section implements an unregistered operation.
// 
wire local_bb2_or296_i_valid_out;
wire local_bb2_or296_i_stall_in;
 reg local_bb2_or296_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u128_valid_out;
wire local_bb2_var__u128_stall_in;
 reg local_bb2_var__u128_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i721_valid_out;
wire local_bb2_lor_ext_i721_stall_in;
 reg local_bb2_lor_ext_i721_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i723_valid_out;
wire local_bb2_reduction_0_i723_stall_in;
 reg local_bb2_reduction_0_i723_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i721_inputs_ready;
wire local_bb2_lor_ext_i721_stall_local;
wire [31:0] local_bb2_lor_ext_i721;

assign local_bb2_lor_ext_i721_inputs_ready = (rnode_175to176_bb2_and35_i652_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_not_cmp38_i_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_and270_i718_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_add246_i_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_var__u107_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2__26_i665_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2__26_i665_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_cmp227_i_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_not__46_i716_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_shr272_i_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2__26_i665_0_valid_out_2_NO_SHIFT_REG & rnode_175to176_bb2_cmp227_i_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2_cmp297_i_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_cmp300_i_0_valid_out_NO_SHIFT_REG);
assign local_bb2_lor_ext_i721 = (local_bb2_cmp29749_i | local_bb2_and303_i);
assign local_bb2_or296_i_valid_out = 1'b1;
assign local_bb2_var__u128_valid_out = 1'b1;
assign local_bb2_lor_ext_i721_valid_out = 1'b1;
assign local_bb2_reduction_0_i723_valid_out = 1'b1;
assign rnode_175to176_bb2_and35_i652_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not_cmp38_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and270_i718_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add246_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u107_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i665_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i665_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp227_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not__46_i716_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_shr272_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i665_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp227_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp297_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp300_i_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_or296_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u128_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_lor_ext_i721_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i723_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_or296_i_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i721_inputs_ready & (local_bb2_or296_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_or296_i_stall_in)) & local_bb2_lor_ext_i721_stall_local);
		local_bb2_var__u128_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i721_inputs_ready & (local_bb2_var__u128_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u128_stall_in)) & local_bb2_lor_ext_i721_stall_local);
		local_bb2_lor_ext_i721_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i721_inputs_ready & (local_bb2_lor_ext_i721_consumed_0_NO_SHIFT_REG | ~(local_bb2_lor_ext_i721_stall_in)) & local_bb2_lor_ext_i721_stall_local);
		local_bb2_reduction_0_i723_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i721_inputs_ready & (local_bb2_reduction_0_i723_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i723_stall_in)) & local_bb2_lor_ext_i721_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_or296_i1809_valid_out;
wire local_bb2_or296_i1809_stall_in;
 reg local_bb2_or296_i1809_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u131_valid_out;
wire local_bb2_var__u131_stall_in;
 reg local_bb2_var__u131_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i1815_valid_out;
wire local_bb2_lor_ext_i1815_stall_in;
 reg local_bb2_lor_ext_i1815_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i1819_valid_out;
wire local_bb2_reduction_0_i1819_stall_in;
 reg local_bb2_reduction_0_i1819_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i1815_inputs_ready;
wire local_bb2_lor_ext_i1815_stall_local;
wire [31:0] local_bb2_lor_ext_i1815;

assign local_bb2_lor_ext_i1815_inputs_ready = (rnode_175to176_bb2_and35_i1664_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_not_cmp38_i1772_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_and270_i1798_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_add246_i1784_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_var__u102_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2__26_i1679_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2__26_i1679_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_add246_i1784_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2_notrhs_i1789_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_cmp227_i1778_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_shr272_i1796_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2__26_i1679_0_valid_out_2_NO_SHIFT_REG & rnode_175to176_bb2_cmp227_i1778_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2_cmp297_i1810_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_cmp300_i1811_0_valid_out_NO_SHIFT_REG);
assign local_bb2_lor_ext_i1815 = (local_bb2_cmp29749_i1814 | local_bb2_and303_i1813);
assign local_bb2_or296_i1809_valid_out = 1'b1;
assign local_bb2_var__u131_valid_out = 1'b1;
assign local_bb2_lor_ext_i1815_valid_out = 1'b1;
assign local_bb2_reduction_0_i1819_valid_out = 1'b1;
assign rnode_175to176_bb2_and35_i1664_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not_cmp38_i1772_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and270_i1798_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add246_i1784_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u102_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1679_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1679_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add246_i1784_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_notrhs_i1789_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp227_i1778_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_shr272_i1796_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1679_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp227_i1778_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp297_i1810_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp300_i1811_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_or296_i1809_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u131_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_lor_ext_i1815_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i1819_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_or296_i1809_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1815_inputs_ready & (local_bb2_or296_i1809_consumed_0_NO_SHIFT_REG | ~(local_bb2_or296_i1809_stall_in)) & local_bb2_lor_ext_i1815_stall_local);
		local_bb2_var__u131_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1815_inputs_ready & (local_bb2_var__u131_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u131_stall_in)) & local_bb2_lor_ext_i1815_stall_local);
		local_bb2_lor_ext_i1815_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1815_inputs_ready & (local_bb2_lor_ext_i1815_consumed_0_NO_SHIFT_REG | ~(local_bb2_lor_ext_i1815_stall_in)) & local_bb2_lor_ext_i1815_stall_local);
		local_bb2_reduction_0_i1819_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1815_inputs_ready & (local_bb2_reduction_0_i1819_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i1819_stall_in)) & local_bb2_lor_ext_i1815_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_or295_i1260_stall_local;
wire [31:0] local_bb2_or295_i1260;

assign local_bb2_or295_i1260 = (local_bb2_or294_i1259 | local_bb2_and293_i1258);

// This section implements an unregistered operation.
// 
wire local_bb2_and302_i1264_stall_local;
wire [31:0] local_bb2_and302_i1264;

assign local_bb2_and302_i1264 = (local_bb2_conv300_i1263 & local_bb2_and293_i1258);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i248_stall_local;
wire [31:0] local_bb2_or295_i248;

assign local_bb2_or295_i248 = (local_bb2_or294_i247 | local_bb2_and293_i246);

// This section implements an unregistered operation.
// 
wire local_bb2_and302_i252_stall_local;
wire [31:0] local_bb2_and302_i252;

assign local_bb2_and302_i252 = (local_bb2_conv300_i251 & local_bb2_and293_i246);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_or296_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_or296_i_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_or296_i_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_or296_i_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_or296_i_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_or296_i_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_or296_i_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_or296_i_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_or296_i),
	.data_out(rnode_176to177_bb2_or296_i_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_or296_i_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_or296_i_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_or296_i_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_or296_i_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_or296_i_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or296_i_stall_in = 1'b0;
assign rnode_176to177_bb2_or296_i_0_NO_SHIFT_REG = rnode_176to177_bb2_or296_i_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_or296_i_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_or296_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_var__u128_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u128_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_var__u128_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u128_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_var__u128_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u128_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u128_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u128_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_var__u128_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_var__u128_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_var__u128_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_var__u128_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_var__u128_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_var__u128),
	.data_out(rnode_176to177_bb2_var__u128_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_var__u128_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_var__u128_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_var__u128_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_var__u128_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_var__u128_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u128_stall_in = 1'b0;
assign rnode_176to177_bb2_var__u128_0_NO_SHIFT_REG = rnode_176to177_bb2_var__u128_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_var__u128_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_var__u128_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_lor_ext_i721_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i721_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_lor_ext_i721_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i721_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_lor_ext_i721_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i721_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i721_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i721_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_lor_ext_i721_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_lor_ext_i721_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_lor_ext_i721_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_lor_ext_i721_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_lor_ext_i721_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_lor_ext_i721),
	.data_out(rnode_176to177_bb2_lor_ext_i721_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_lor_ext_i721_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_lor_ext_i721_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_lor_ext_i721_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_lor_ext_i721_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_lor_ext_i721_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lor_ext_i721_stall_in = 1'b0;
assign rnode_176to177_bb2_lor_ext_i721_0_NO_SHIFT_REG = rnode_176to177_bb2_lor_ext_i721_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_lor_ext_i721_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_lor_ext_i721_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_reduction_0_i723_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i723_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_reduction_0_i723_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i723_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_reduction_0_i723_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i723_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i723_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i723_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_reduction_0_i723_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_reduction_0_i723_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_reduction_0_i723_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_reduction_0_i723_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_reduction_0_i723_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i723),
	.data_out(rnode_176to177_bb2_reduction_0_i723_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_reduction_0_i723_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_reduction_0_i723_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_reduction_0_i723_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_reduction_0_i723_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_reduction_0_i723_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i723_stall_in = 1'b0;
assign rnode_176to177_bb2_reduction_0_i723_0_NO_SHIFT_REG = rnode_176to177_bb2_reduction_0_i723_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_reduction_0_i723_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_reduction_0_i723_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_or296_i1809_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i1809_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_or296_i1809_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i1809_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_or296_i1809_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i1809_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i1809_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or296_i1809_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_or296_i1809_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_or296_i1809_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_or296_i1809_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_or296_i1809_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_or296_i1809_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_or296_i1809),
	.data_out(rnode_176to177_bb2_or296_i1809_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_or296_i1809_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_or296_i1809_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_or296_i1809_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_or296_i1809_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_or296_i1809_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or296_i1809_stall_in = 1'b0;
assign rnode_176to177_bb2_or296_i1809_0_NO_SHIFT_REG = rnode_176to177_bb2_or296_i1809_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_or296_i1809_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_or296_i1809_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_var__u131_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u131_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_var__u131_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u131_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_var__u131_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u131_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u131_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u131_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_var__u131_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_var__u131_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_var__u131_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_var__u131_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_var__u131_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_var__u131),
	.data_out(rnode_176to177_bb2_var__u131_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_var__u131_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_var__u131_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_var__u131_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_var__u131_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_var__u131_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u131_stall_in = 1'b0;
assign rnode_176to177_bb2_var__u131_0_NO_SHIFT_REG = rnode_176to177_bb2_var__u131_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_var__u131_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_var__u131_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_lor_ext_i1815_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1815_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_lor_ext_i1815_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1815_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_lor_ext_i1815_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1815_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1815_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1815_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_lor_ext_i1815_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_lor_ext_i1815_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_lor_ext_i1815_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_lor_ext_i1815_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_lor_ext_i1815_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_lor_ext_i1815),
	.data_out(rnode_176to177_bb2_lor_ext_i1815_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_lor_ext_i1815_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_lor_ext_i1815_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_lor_ext_i1815_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_lor_ext_i1815_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_lor_ext_i1815_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lor_ext_i1815_stall_in = 1'b0;
assign rnode_176to177_bb2_lor_ext_i1815_0_NO_SHIFT_REG = rnode_176to177_bb2_lor_ext_i1815_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_lor_ext_i1815_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_lor_ext_i1815_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_reduction_0_i1819_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1819_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_reduction_0_i1819_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1819_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_reduction_0_i1819_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1819_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1819_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1819_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_reduction_0_i1819_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_reduction_0_i1819_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_reduction_0_i1819_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_reduction_0_i1819_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_reduction_0_i1819_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i1819),
	.data_out(rnode_176to177_bb2_reduction_0_i1819_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_reduction_0_i1819_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_reduction_0_i1819_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_reduction_0_i1819_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_reduction_0_i1819_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_reduction_0_i1819_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i1819_stall_in = 1'b0;
assign rnode_176to177_bb2_reduction_0_i1819_0_NO_SHIFT_REG = rnode_176to177_bb2_reduction_0_i1819_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_reduction_0_i1819_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_reduction_0_i1819_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i1260_valid_out;
wire local_bb2_or295_i1260_stall_in;
 reg local_bb2_or295_i1260_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u134_valid_out;
wire local_bb2_var__u134_stall_in;
 reg local_bb2_var__u134_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i1266_valid_out;
wire local_bb2_lor_ext_i1266_stall_in;
 reg local_bb2_lor_ext_i1266_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i1270_valid_out;
wire local_bb2_reduction_0_i1270_stall_in;
 reg local_bb2_reduction_0_i1270_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i1266_inputs_ready;
wire local_bb2_lor_ext_i1266_stall_local;
wire [31:0] local_bb2_lor_ext_i1266;

assign local_bb2_lor_ext_i1266_inputs_ready = (rnode_175to176_bb2_and35_i1115_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_not_cmp37_i1223_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_and269_i1249_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_add245_i1235_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_var__u111_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2__26_i1130_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2__26_i1130_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_add245_i1235_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2_notrhs_i1240_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_cmp226_i1229_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_shr271_i1247_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2__26_i1130_0_valid_out_2_NO_SHIFT_REG & rnode_175to176_bb2_cmp226_i1229_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2_cmp296_i1261_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_cmp299_i1262_0_valid_out_NO_SHIFT_REG);
assign local_bb2_lor_ext_i1266 = (local_bb2_cmp29649_i1265 | local_bb2_and302_i1264);
assign local_bb2_or295_i1260_valid_out = 1'b1;
assign local_bb2_var__u134_valid_out = 1'b1;
assign local_bb2_lor_ext_i1266_valid_out = 1'b1;
assign local_bb2_reduction_0_i1270_valid_out = 1'b1;
assign rnode_175to176_bb2_and35_i1115_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not_cmp37_i1223_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and269_i1249_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add245_i1235_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u111_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1130_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1130_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add245_i1235_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_notrhs_i1240_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp226_i1229_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_shr271_i1247_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i1130_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp226_i1229_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp296_i1261_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp299_i1262_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_or295_i1260_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u134_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_lor_ext_i1266_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i1270_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_or295_i1260_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1266_inputs_ready & (local_bb2_or295_i1260_consumed_0_NO_SHIFT_REG | ~(local_bb2_or295_i1260_stall_in)) & local_bb2_lor_ext_i1266_stall_local);
		local_bb2_var__u134_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1266_inputs_ready & (local_bb2_var__u134_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u134_stall_in)) & local_bb2_lor_ext_i1266_stall_local);
		local_bb2_lor_ext_i1266_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1266_inputs_ready & (local_bb2_lor_ext_i1266_consumed_0_NO_SHIFT_REG | ~(local_bb2_lor_ext_i1266_stall_in)) & local_bb2_lor_ext_i1266_stall_local);
		local_bb2_reduction_0_i1270_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1266_inputs_ready & (local_bb2_reduction_0_i1270_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i1270_stall_in)) & local_bb2_lor_ext_i1266_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_or295_i248_valid_out;
wire local_bb2_or295_i248_stall_in;
 reg local_bb2_or295_i248_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u135_valid_out;
wire local_bb2_var__u135_stall_in;
 reg local_bb2_var__u135_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i254_valid_out;
wire local_bb2_lor_ext_i254_stall_in;
 reg local_bb2_lor_ext_i254_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i258_valid_out;
wire local_bb2_reduction_0_i258_stall_in;
 reg local_bb2_reduction_0_i258_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i254_inputs_ready;
wire local_bb2_lor_ext_i254_stall_local;
wire [31:0] local_bb2_lor_ext_i254;

assign local_bb2_lor_ext_i254_inputs_ready = (rnode_175to176_bb2_and35_i103_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_not_cmp37_i211_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_and269_i237_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_add245_i223_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_var__u114_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2__26_i118_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2__26_i118_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_add245_i223_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2_notrhs_i228_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_cmp226_i217_0_valid_out_1_NO_SHIFT_REG & rnode_175to176_bb2_shr271_i235_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2__26_i118_0_valid_out_2_NO_SHIFT_REG & rnode_175to176_bb2_cmp226_i217_0_valid_out_0_NO_SHIFT_REG & rnode_175to176_bb2_cmp296_i249_0_valid_out_NO_SHIFT_REG & rnode_175to176_bb2_cmp299_i250_0_valid_out_NO_SHIFT_REG);
assign local_bb2_lor_ext_i254 = (local_bb2_cmp29649_i253 | local_bb2_and302_i252);
assign local_bb2_or295_i248_valid_out = 1'b1;
assign local_bb2_var__u135_valid_out = 1'b1;
assign local_bb2_lor_ext_i254_valid_out = 1'b1;
assign local_bb2_reduction_0_i258_valid_out = 1'b1;
assign rnode_175to176_bb2_and35_i103_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_not_cmp37_i211_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_and269_i237_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add245_i223_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_var__u114_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i118_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i118_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_add245_i223_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_notrhs_i228_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp226_i217_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_shr271_i235_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2__26_i118_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp226_i217_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp296_i249_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_175to176_bb2_cmp299_i250_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_or295_i248_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u135_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_lor_ext_i254_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i258_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_or295_i248_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i254_inputs_ready & (local_bb2_or295_i248_consumed_0_NO_SHIFT_REG | ~(local_bb2_or295_i248_stall_in)) & local_bb2_lor_ext_i254_stall_local);
		local_bb2_var__u135_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i254_inputs_ready & (local_bb2_var__u135_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u135_stall_in)) & local_bb2_lor_ext_i254_stall_local);
		local_bb2_lor_ext_i254_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i254_inputs_ready & (local_bb2_lor_ext_i254_consumed_0_NO_SHIFT_REG | ~(local_bb2_lor_ext_i254_stall_in)) & local_bb2_lor_ext_i254_stall_local);
		local_bb2_reduction_0_i258_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i254_inputs_ready & (local_bb2_reduction_0_i258_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i258_stall_in)) & local_bb2_lor_ext_i254_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext315_i_stall_local;
wire [31:0] local_bb2_lnot_ext315_i;

assign local_bb2_lnot_ext315_i = (rnode_176to177_bb2_var__u128_0_NO_SHIFT_REG ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext315_i1818_stall_local;
wire [31:0] local_bb2_lnot_ext315_i1818;

assign local_bb2_lnot_ext315_i1818 = (rnode_176to177_bb2_var__u131_0_NO_SHIFT_REG ^ 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_or295_i1260_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i1260_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_or295_i1260_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i1260_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_or295_i1260_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i1260_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i1260_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i1260_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_or295_i1260_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_or295_i1260_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_or295_i1260_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_or295_i1260_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_or295_i1260_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_or295_i1260),
	.data_out(rnode_176to177_bb2_or295_i1260_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_or295_i1260_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_or295_i1260_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_or295_i1260_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_or295_i1260_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_or295_i1260_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or295_i1260_stall_in = 1'b0;
assign rnode_176to177_bb2_or295_i1260_0_NO_SHIFT_REG = rnode_176to177_bb2_or295_i1260_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_or295_i1260_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_or295_i1260_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_var__u134_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u134_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_var__u134_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u134_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_var__u134_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u134_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u134_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u134_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_var__u134_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_var__u134_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_var__u134_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_var__u134_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_var__u134_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_var__u134),
	.data_out(rnode_176to177_bb2_var__u134_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_var__u134_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_var__u134_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_var__u134_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_var__u134_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_var__u134_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u134_stall_in = 1'b0;
assign rnode_176to177_bb2_var__u134_0_NO_SHIFT_REG = rnode_176to177_bb2_var__u134_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_var__u134_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_var__u134_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_lor_ext_i1266_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1266_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_lor_ext_i1266_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1266_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_lor_ext_i1266_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1266_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1266_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i1266_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_lor_ext_i1266_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_lor_ext_i1266_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_lor_ext_i1266_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_lor_ext_i1266_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_lor_ext_i1266_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_lor_ext_i1266),
	.data_out(rnode_176to177_bb2_lor_ext_i1266_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_lor_ext_i1266_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_lor_ext_i1266_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_lor_ext_i1266_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_lor_ext_i1266_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_lor_ext_i1266_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lor_ext_i1266_stall_in = 1'b0;
assign rnode_176to177_bb2_lor_ext_i1266_0_NO_SHIFT_REG = rnode_176to177_bb2_lor_ext_i1266_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_lor_ext_i1266_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_lor_ext_i1266_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_reduction_0_i1270_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1270_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_reduction_0_i1270_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1270_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_reduction_0_i1270_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1270_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1270_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i1270_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_reduction_0_i1270_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_reduction_0_i1270_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_reduction_0_i1270_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_reduction_0_i1270_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_reduction_0_i1270_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i1270),
	.data_out(rnode_176to177_bb2_reduction_0_i1270_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_reduction_0_i1270_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_reduction_0_i1270_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_reduction_0_i1270_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_reduction_0_i1270_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_reduction_0_i1270_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i1270_stall_in = 1'b0;
assign rnode_176to177_bb2_reduction_0_i1270_0_NO_SHIFT_REG = rnode_176to177_bb2_reduction_0_i1270_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_reduction_0_i1270_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_reduction_0_i1270_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_or295_i248_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i248_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_or295_i248_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i248_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_or295_i248_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i248_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i248_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_or295_i248_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_or295_i248_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_or295_i248_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_or295_i248_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_or295_i248_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_or295_i248_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_or295_i248),
	.data_out(rnode_176to177_bb2_or295_i248_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_or295_i248_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_or295_i248_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_or295_i248_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_or295_i248_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_or295_i248_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or295_i248_stall_in = 1'b0;
assign rnode_176to177_bb2_or295_i248_0_NO_SHIFT_REG = rnode_176to177_bb2_or295_i248_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_or295_i248_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_or295_i248_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_var__u135_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u135_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_var__u135_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u135_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_var__u135_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u135_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u135_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_var__u135_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_var__u135_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_var__u135_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_var__u135_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_var__u135_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_var__u135_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_var__u135),
	.data_out(rnode_176to177_bb2_var__u135_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_var__u135_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_var__u135_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_var__u135_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_var__u135_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_var__u135_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u135_stall_in = 1'b0;
assign rnode_176to177_bb2_var__u135_0_NO_SHIFT_REG = rnode_176to177_bb2_var__u135_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_var__u135_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_var__u135_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_lor_ext_i254_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i254_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_lor_ext_i254_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i254_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_lor_ext_i254_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i254_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i254_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_lor_ext_i254_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_lor_ext_i254_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_lor_ext_i254_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_lor_ext_i254_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_lor_ext_i254_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_lor_ext_i254_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_lor_ext_i254),
	.data_out(rnode_176to177_bb2_lor_ext_i254_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_lor_ext_i254_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_lor_ext_i254_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_lor_ext_i254_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_lor_ext_i254_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_lor_ext_i254_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lor_ext_i254_stall_in = 1'b0;
assign rnode_176to177_bb2_lor_ext_i254_0_NO_SHIFT_REG = rnode_176to177_bb2_lor_ext_i254_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_lor_ext_i254_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_lor_ext_i254_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_176to177_bb2_reduction_0_i258_0_valid_out_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i258_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_reduction_0_i258_0_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i258_0_reg_177_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_176to177_bb2_reduction_0_i258_0_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i258_0_valid_out_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i258_0_stall_in_reg_177_NO_SHIFT_REG;
 logic rnode_176to177_bb2_reduction_0_i258_0_stall_out_reg_177_NO_SHIFT_REG;

acl_data_fifo rnode_176to177_bb2_reduction_0_i258_0_reg_177_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_176to177_bb2_reduction_0_i258_0_reg_177_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_176to177_bb2_reduction_0_i258_0_stall_in_reg_177_NO_SHIFT_REG),
	.valid_out(rnode_176to177_bb2_reduction_0_i258_0_valid_out_reg_177_NO_SHIFT_REG),
	.stall_out(rnode_176to177_bb2_reduction_0_i258_0_stall_out_reg_177_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i258),
	.data_out(rnode_176to177_bb2_reduction_0_i258_0_reg_177_NO_SHIFT_REG)
);

defparam rnode_176to177_bb2_reduction_0_i258_0_reg_177_fifo.DEPTH = 1;
defparam rnode_176to177_bb2_reduction_0_i258_0_reg_177_fifo.DATA_WIDTH = 32;
defparam rnode_176to177_bb2_reduction_0_i258_0_reg_177_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_176to177_bb2_reduction_0_i258_0_reg_177_fifo.IMPL = "shift_reg";

assign rnode_176to177_bb2_reduction_0_i258_0_reg_177_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i258_stall_in = 1'b0;
assign rnode_176to177_bb2_reduction_0_i258_0_NO_SHIFT_REG = rnode_176to177_bb2_reduction_0_i258_0_reg_177_NO_SHIFT_REG;
assign rnode_176to177_bb2_reduction_0_i258_0_stall_in_reg_177_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_reduction_0_i258_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_1_i724_stall_local;
wire [31:0] local_bb2_reduction_1_i724;

assign local_bb2_reduction_1_i724 = (local_bb2_lnot_ext315_i & rnode_176to177_bb2_lor_ext_i721_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_1_i1820_stall_local;
wire [31:0] local_bb2_reduction_1_i1820;

assign local_bb2_reduction_1_i1820 = (local_bb2_lnot_ext315_i1818 & rnode_176to177_bb2_lor_ext_i1815_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext314_i1269_stall_local;
wire [31:0] local_bb2_lnot_ext314_i1269;

assign local_bb2_lnot_ext314_i1269 = (rnode_176to177_bb2_var__u134_0_NO_SHIFT_REG ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext314_i257_stall_local;
wire [31:0] local_bb2_lnot_ext314_i257;

assign local_bb2_lnot_ext314_i257 = (rnode_176to177_bb2_var__u135_0_NO_SHIFT_REG ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i725_stall_local;
wire [31:0] local_bb2_reduction_2_i725;

assign local_bb2_reduction_2_i725 = (rnode_176to177_bb2_reduction_0_i723_0_NO_SHIFT_REG & local_bb2_reduction_1_i724);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i1821_stall_local;
wire [31:0] local_bb2_reduction_2_i1821;

assign local_bb2_reduction_2_i1821 = (rnode_176to177_bb2_reduction_0_i1819_0_NO_SHIFT_REG & local_bb2_reduction_1_i1820);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_1_i1271_stall_local;
wire [31:0] local_bb2_reduction_1_i1271;

assign local_bb2_reduction_1_i1271 = (local_bb2_lnot_ext314_i1269 & rnode_176to177_bb2_lor_ext_i1266_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_1_i259_stall_local;
wire [31:0] local_bb2_reduction_1_i259;

assign local_bb2_reduction_1_i259 = (local_bb2_lnot_ext314_i257 & rnode_176to177_bb2_lor_ext_i254_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_add321_i_valid_out;
wire local_bb2_add321_i_stall_in;
wire local_bb2_add321_i_inputs_ready;
wire local_bb2_add321_i_stall_local;
wire [31:0] local_bb2_add321_i;

assign local_bb2_add321_i_inputs_ready = (rnode_176to177_bb2_or296_i_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_reduction_0_i723_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_var__u128_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_lor_ext_i721_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add321_i = (local_bb2_reduction_2_i725 + rnode_176to177_bb2_or296_i_0_NO_SHIFT_REG);
assign local_bb2_add321_i_valid_out = 1'b1;
assign rnode_176to177_bb2_or296_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_reduction_0_i723_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_var__u128_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_lor_ext_i721_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_add321_i1822_valid_out;
wire local_bb2_add321_i1822_stall_in;
wire local_bb2_add321_i1822_inputs_ready;
wire local_bb2_add321_i1822_stall_local;
wire [31:0] local_bb2_add321_i1822;

assign local_bb2_add321_i1822_inputs_ready = (rnode_176to177_bb2_or296_i1809_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_reduction_0_i1819_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_var__u131_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_lor_ext_i1815_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add321_i1822 = (local_bb2_reduction_2_i1821 + rnode_176to177_bb2_or296_i1809_0_NO_SHIFT_REG);
assign local_bb2_add321_i1822_valid_out = 1'b1;
assign rnode_176to177_bb2_or296_i1809_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_reduction_0_i1819_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_var__u131_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_lor_ext_i1815_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i1272_stall_local;
wire [31:0] local_bb2_reduction_2_i1272;

assign local_bb2_reduction_2_i1272 = (rnode_176to177_bb2_reduction_0_i1270_0_NO_SHIFT_REG & local_bb2_reduction_1_i1271);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i260_stall_local;
wire [31:0] local_bb2_reduction_2_i260;

assign local_bb2_reduction_2_i260 = (rnode_176to177_bb2_reduction_0_i258_0_NO_SHIFT_REG & local_bb2_reduction_1_i259);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb2_add321_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add321_i_0_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add321_i_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb2_add321_i_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb2_add321_i_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb2_add321_i_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb2_add321_i_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb2_add321_i_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb2_add321_i),
	.data_out(rnode_177to178_bb2_add321_i_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb2_add321_i_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb2_add321_i_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb2_add321_i_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb2_add321_i_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb2_add321_i_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add321_i_stall_in = 1'b0;
assign rnode_177to178_bb2_add321_i_0_NO_SHIFT_REG = rnode_177to178_bb2_add321_i_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_add321_i_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add321_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb2_add321_i1822_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add321_i1822_0_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add321_i1822_1_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add321_i1822_2_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add321_i1822_3_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add321_i1822_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add321_i1822_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb2_add321_i1822_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb2_add321_i1822_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb2_add321_i1822_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb2_add321_i1822_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb2_add321_i1822_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb2_add321_i1822),
	.data_out(rnode_177to178_bb2_add321_i1822_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb2_add321_i1822_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb2_add321_i1822_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb2_add321_i1822_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb2_add321_i1822_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb2_add321_i1822_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add321_i1822_stall_in = 1'b0;
assign rnode_177to178_bb2_add321_i1822_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add321_i1822_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add321_i1822_0_NO_SHIFT_REG = rnode_177to178_bb2_add321_i1822_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_add321_i1822_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add321_i1822_1_NO_SHIFT_REG = rnode_177to178_bb2_add321_i1822_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_add321_i1822_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add321_i1822_2_NO_SHIFT_REG = rnode_177to178_bb2_add321_i1822_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_add321_i1822_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add321_i1822_3_NO_SHIFT_REG = rnode_177to178_bb2_add321_i1822_0_reg_178_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_add320_i1273_valid_out;
wire local_bb2_add320_i1273_stall_in;
wire local_bb2_add320_i1273_inputs_ready;
wire local_bb2_add320_i1273_stall_local;
wire [31:0] local_bb2_add320_i1273;

assign local_bb2_add320_i1273_inputs_ready = (rnode_176to177_bb2_or295_i1260_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_reduction_0_i1270_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_var__u134_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_lor_ext_i1266_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add320_i1273 = (local_bb2_reduction_2_i1272 + rnode_176to177_bb2_or295_i1260_0_NO_SHIFT_REG);
assign local_bb2_add320_i1273_valid_out = 1'b1;
assign rnode_176to177_bb2_or295_i1260_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_reduction_0_i1270_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_var__u134_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_lor_ext_i1266_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_add320_i261_valid_out;
wire local_bb2_add320_i261_stall_in;
wire local_bb2_add320_i261_inputs_ready;
wire local_bb2_add320_i261_stall_local;
wire [31:0] local_bb2_add320_i261;

assign local_bb2_add320_i261_inputs_ready = (rnode_176to177_bb2_or295_i248_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_reduction_0_i258_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_var__u135_0_valid_out_NO_SHIFT_REG & rnode_176to177_bb2_lor_ext_i254_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add320_i261 = (local_bb2_reduction_2_i260 + rnode_176to177_bb2_or295_i248_0_NO_SHIFT_REG);
assign local_bb2_add320_i261_valid_out = 1'b1;
assign rnode_176to177_bb2_or295_i248_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_reduction_0_i258_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_var__u135_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_176to177_bb2_lor_ext_i254_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_178to184_bb2_add321_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add321_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_178to184_bb2_add321_i_0_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add321_i_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to184_bb2_add321_i_0_reg_184_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add321_i_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add321_i_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add321_i_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_178to184_bb2_add321_i_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to184_bb2_add321_i_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to184_bb2_add321_i_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_178to184_bb2_add321_i_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_178to184_bb2_add321_i_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb2_add321_i_0_NO_SHIFT_REG),
	.data_out(rnode_178to184_bb2_add321_i_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_178to184_bb2_add321_i_0_reg_184_fifo.DEPTH = 6;
defparam rnode_178to184_bb2_add321_i_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_178to184_bb2_add321_i_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to184_bb2_add321_i_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_178to184_bb2_add321_i_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add321_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to184_bb2_add321_i_0_NO_SHIFT_REG = rnode_178to184_bb2_add321_i_0_reg_184_NO_SHIFT_REG;
assign rnode_178to184_bb2_add321_i_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_178to184_bb2_add321_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and_i1458_stall_local;
wire [31:0] local_bb2_and_i1458;

assign local_bb2_and_i1458 = (rnode_177to178_bb2_add321_i1822_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and10_i1464_stall_local;
wire [31:0] local_bb2_and10_i1464;

assign local_bb2_and10_i1464 = (rnode_177to178_bb2_add321_i1822_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb2_add320_i1273_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add320_i1273_0_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add320_i1273_1_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add320_i1273_2_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add320_i1273_3_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add320_i1273_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_valid_out_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_stall_in_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i1273_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb2_add320_i1273_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb2_add320_i1273_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb2_add320_i1273_0_stall_in_0_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb2_add320_i1273_0_valid_out_0_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb2_add320_i1273_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb2_add320_i1273),
	.data_out(rnode_177to178_bb2_add320_i1273_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb2_add320_i1273_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb2_add320_i1273_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb2_add320_i1273_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb2_add320_i1273_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb2_add320_i1273_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add320_i1273_stall_in = 1'b0;
assign rnode_177to178_bb2_add320_i1273_0_stall_in_0_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add320_i1273_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add320_i1273_0_NO_SHIFT_REG = rnode_177to178_bb2_add320_i1273_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_add320_i1273_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add320_i1273_1_NO_SHIFT_REG = rnode_177to178_bb2_add320_i1273_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_add320_i1273_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add320_i1273_2_NO_SHIFT_REG = rnode_177to178_bb2_add320_i1273_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_add320_i1273_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add320_i1273_3_NO_SHIFT_REG = rnode_177to178_bb2_add320_i1273_0_reg_178_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_177to178_bb2_add320_i261_0_valid_out_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i261_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add320_i261_0_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i261_0_reg_178_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_177to178_bb2_add320_i261_0_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i261_0_valid_out_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i261_0_stall_in_reg_178_NO_SHIFT_REG;
 logic rnode_177to178_bb2_add320_i261_0_stall_out_reg_178_NO_SHIFT_REG;

acl_data_fifo rnode_177to178_bb2_add320_i261_0_reg_178_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_177to178_bb2_add320_i261_0_reg_178_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_177to178_bb2_add320_i261_0_stall_in_reg_178_NO_SHIFT_REG),
	.valid_out(rnode_177to178_bb2_add320_i261_0_valid_out_reg_178_NO_SHIFT_REG),
	.stall_out(rnode_177to178_bb2_add320_i261_0_stall_out_reg_178_NO_SHIFT_REG),
	.data_in(local_bb2_add320_i261),
	.data_out(rnode_177to178_bb2_add320_i261_0_reg_178_NO_SHIFT_REG)
);

defparam rnode_177to178_bb2_add320_i261_0_reg_178_fifo.DEPTH = 1;
defparam rnode_177to178_bb2_add320_i261_0_reg_178_fifo.DATA_WIDTH = 32;
defparam rnode_177to178_bb2_add320_i261_0_reg_178_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_177to178_bb2_add320_i261_0_reg_178_fifo.IMPL = "shift_reg";

assign rnode_177to178_bb2_add320_i261_0_reg_178_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add320_i261_stall_in = 1'b0;
assign rnode_177to178_bb2_add320_i261_0_NO_SHIFT_REG = rnode_177to178_bb2_add320_i261_0_reg_178_NO_SHIFT_REG;
assign rnode_177to178_bb2_add320_i261_0_stall_in_reg_178_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add320_i261_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb2_add321_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add321_i_0_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add321_i_1_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add321_i_2_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add321_i_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_valid_out_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_stall_in_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add321_i_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb2_add321_i_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb2_add321_i_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb2_add321_i_0_stall_in_0_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb2_add321_i_0_valid_out_0_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb2_add321_i_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(rnode_178to184_bb2_add321_i_0_NO_SHIFT_REG),
	.data_out(rnode_184to185_bb2_add321_i_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb2_add321_i_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb2_add321_i_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb2_add321_i_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb2_add321_i_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb2_add321_i_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to184_bb2_add321_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add321_i_0_stall_in_0_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add321_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add321_i_0_NO_SHIFT_REG = rnode_184to185_bb2_add321_i_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb2_add321_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add321_i_1_NO_SHIFT_REG = rnode_184to185_bb2_add321_i_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb2_add321_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add321_i_2_NO_SHIFT_REG = rnode_184to185_bb2_add321_i_0_reg_185_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i1459_stall_local;
wire [31:0] local_bb2_shr_i1459;

assign local_bb2_shr_i1459 = (local_bb2_and_i1458 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp13_i1466_stall_local;
wire local_bb2_cmp13_i1466;

assign local_bb2_cmp13_i1466 = (local_bb2_and10_i1464 > local_bb2_and12_i1465);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i910_stall_local;
wire [31:0] local_bb2_and_i910;

assign local_bb2_and_i910 = (rnode_177to178_bb2_add320_i1273_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and10_i916_stall_local;
wire [31:0] local_bb2_and10_i916;

assign local_bb2_and10_i916 = (rnode_177to178_bb2_add320_i1273_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 6
//  * capacity = 6
 logic rnode_178to184_bb2_add320_i261_0_valid_out_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add320_i261_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_178to184_bb2_add320_i261_0_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add320_i261_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to184_bb2_add320_i261_0_reg_184_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add320_i261_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add320_i261_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_178to184_bb2_add320_i261_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_178to184_bb2_add320_i261_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to184_bb2_add320_i261_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to184_bb2_add320_i261_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_178to184_bb2_add320_i261_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_178to184_bb2_add320_i261_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(rnode_177to178_bb2_add320_i261_0_NO_SHIFT_REG),
	.data_out(rnode_178to184_bb2_add320_i261_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_178to184_bb2_add320_i261_0_reg_184_fifo.DEPTH = 6;
defparam rnode_178to184_bb2_add320_i261_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_178to184_bb2_add320_i261_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to184_bb2_add320_i261_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_178to184_bb2_add320_i261_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_177to178_bb2_add320_i261_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_178to184_bb2_add320_i261_0_NO_SHIFT_REG = rnode_178to184_bb2_add320_i261_0_reg_184_NO_SHIFT_REG;
assign rnode_178to184_bb2_add320_i261_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_178to184_bb2_add320_i261_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and_i446_stall_local;
wire [31:0] local_bb2_and_i446;

assign local_bb2_and_i446 = (rnode_184to185_bb2_add321_i_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and10_i452_stall_local;
wire [31:0] local_bb2_and10_i452;

assign local_bb2_and10_i452 = (rnode_184to185_bb2_add321_i_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb2_add321_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add321_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add321_i_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add321_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add321_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add321_i_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add321_i_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add321_i_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add321_i_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add321_i_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add321_i_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb2_add321_i_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb2_add321_i_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb2_add321_i_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb2_add321_i_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb2_add321_i_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_184to185_bb2_add321_i_2_NO_SHIFT_REG),
	.data_out(rnode_185to186_bb2_add321_i_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb2_add321_i_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb2_add321_i_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_185to186_bb2_add321_i_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb2_add321_i_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb2_add321_i_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add321_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add321_i_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add321_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add321_i_0_NO_SHIFT_REG = rnode_185to186_bb2_add321_i_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb2_add321_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add321_i_1_NO_SHIFT_REG = rnode_185to186_bb2_add321_i_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i1462_stall_local;
wire local_bb2_cmp_i1462;

assign local_bb2_cmp_i1462 = (local_bb2_shr_i1459 > local_bb2_shr3_i1461);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp8_i1463_stall_local;
wire local_bb2_cmp8_i1463;

assign local_bb2_cmp8_i1463 = (local_bb2_shr_i1459 == local_bb2_shr3_i1461);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i911_stall_local;
wire [31:0] local_bb2_shr_i911;

assign local_bb2_shr_i911 = (local_bb2_and_i910 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp13_i918_stall_local;
wire local_bb2_cmp13_i918;

assign local_bb2_cmp13_i918 = (local_bb2_and10_i916 > local_bb2_and12_i917);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb2_add320_i261_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i261_0_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i261_1_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i261_2_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i261_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_valid_out_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_stall_in_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i261_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb2_add320_i261_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb2_add320_i261_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb2_add320_i261_0_stall_in_0_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb2_add320_i261_0_valid_out_0_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb2_add320_i261_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(rnode_178to184_bb2_add320_i261_0_NO_SHIFT_REG),
	.data_out(rnode_184to185_bb2_add320_i261_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb2_add320_i261_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb2_add320_i261_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb2_add320_i261_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb2_add320_i261_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb2_add320_i261_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to184_bb2_add320_i261_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add320_i261_0_stall_in_0_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add320_i261_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i261_0_NO_SHIFT_REG = rnode_184to185_bb2_add320_i261_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb2_add320_i261_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i261_1_NO_SHIFT_REG = rnode_184to185_bb2_add320_i261_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb2_add320_i261_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i261_2_NO_SHIFT_REG = rnode_184to185_bb2_add320_i261_0_reg_185_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i447_stall_local;
wire [31:0] local_bb2_shr_i447;

assign local_bb2_shr_i447 = (local_bb2_and_i446 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2___i1467_stall_local;
wire local_bb2___i1467;

assign local_bb2___i1467 = (local_bb2_cmp8_i1463 & local_bb2_cmp13_i1466);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i914_stall_local;
wire local_bb2_cmp_i914;

assign local_bb2_cmp_i914 = (local_bb2_shr_i911 > local_bb2_shr3_i913);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp8_i915_stall_local;
wire local_bb2_cmp8_i915;

assign local_bb2_cmp8_i915 = (local_bb2_shr_i911 == local_bb2_shr3_i913);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i50_stall_local;
wire [31:0] local_bb2_and_i50;

assign local_bb2_and_i50 = (rnode_184to185_bb2_add320_i261_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and10_i_stall_local;
wire [31:0] local_bb2_and10_i;

assign local_bb2_and10_i = (rnode_184to185_bb2_add320_i261_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb2_add320_i261_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i261_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i261_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i261_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i261_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i261_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i261_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i261_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i261_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i261_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i261_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb2_add320_i261_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb2_add320_i261_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb2_add320_i261_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb2_add320_i261_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb2_add320_i261_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_184to185_bb2_add320_i261_2_NO_SHIFT_REG),
	.data_out(rnode_185to186_bb2_add320_i261_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb2_add320_i261_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb2_add320_i261_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_185to186_bb2_add320_i261_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb2_add320_i261_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb2_add320_i261_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i261_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i261_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i261_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i261_0_NO_SHIFT_REG = rnode_185to186_bb2_add320_i261_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb2_add320_i261_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i261_1_NO_SHIFT_REG = rnode_185to186_bb2_add320_i261_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__21_i1468_stall_local;
wire local_bb2__21_i1468;

assign local_bb2__21_i1468 = (local_bb2_cmp_i1462 | local_bb2___i1467);

// This section implements an unregistered operation.
// 
wire local_bb2___i919_stall_local;
wire local_bb2___i919;

assign local_bb2___i919 = (local_bb2_cmp8_i915 & local_bb2_cmp13_i918);

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i51_stall_local;
wire [31:0] local_bb2_shr_i51;

assign local_bb2_shr_i51 = (local_bb2_and_i50 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i1469_stall_local;
wire [31:0] local_bb2__22_i1469;

assign local_bb2__22_i1469 = (local_bb2__21_i1468 ? local_bb2_var__u24 : rnode_177to178_bb2_add321_i1822_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i1469_valid_out;
wire local_bb2__22_i1469_stall_in;
 reg local_bb2__22_i1469_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i1470_valid_out;
wire local_bb2__23_i1470_stall_in;
 reg local_bb2__23_i1470_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i1470_inputs_ready;
wire local_bb2__23_i1470_stall_local;
wire [31:0] local_bb2__23_i1470;

assign local_bb2__23_i1470_inputs_ready = (rnode_177to178_bb2_c0_ene5_0_valid_out_NO_SHIFT_REG & rnode_177to178_bb2_add321_i1822_0_valid_out_2_NO_SHIFT_REG & rnode_177to178_bb2_add321_i1822_0_valid_out_3_NO_SHIFT_REG & rnode_177to178_bb2_add321_i1822_0_valid_out_1_NO_SHIFT_REG & rnode_177to178_bb2_add321_i1822_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2__23_i1470 = (local_bb2__21_i1468 ? rnode_177to178_bb2_add321_i1822_3_NO_SHIFT_REG : local_bb2_var__u24);
assign local_bb2__22_i1469_valid_out = 1'b1;
assign local_bb2__23_i1470_valid_out = 1'b1;
assign rnode_177to178_bb2_c0_ene5_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add321_i1822_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add321_i1822_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add321_i1822_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add321_i1822_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__22_i1469_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__23_i1470_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__22_i1469_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i1470_inputs_ready & (local_bb2__22_i1469_consumed_0_NO_SHIFT_REG | ~(local_bb2__22_i1469_stall_in)) & local_bb2__23_i1470_stall_local);
		local_bb2__23_i1470_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i1470_inputs_ready & (local_bb2__23_i1470_consumed_0_NO_SHIFT_REG | ~(local_bb2__23_i1470_stall_in)) & local_bb2__23_i1470_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2__21_i920_stall_local;
wire local_bb2__21_i920;

assign local_bb2__21_i920 = (local_bb2_cmp_i914 | local_bb2___i919);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb2__22_i1469_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i1469_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__22_i1469_0_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i1469_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i1469_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__22_i1469_1_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i1469_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__22_i1469_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i1469_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i1469_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i1469_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb2__22_i1469_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb2__22_i1469_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb2__22_i1469_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb2__22_i1469_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb2__22_i1469_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb2__22_i1469),
	.data_out(rnode_178to179_bb2__22_i1469_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb2__22_i1469_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb2__22_i1469_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb2__22_i1469_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb2__22_i1469_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb2__22_i1469_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__22_i1469_stall_in = 1'b0;
assign rnode_178to179_bb2__22_i1469_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb2__22_i1469_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__22_i1469_0_NO_SHIFT_REG = rnode_178to179_bb2__22_i1469_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb2__22_i1469_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__22_i1469_1_NO_SHIFT_REG = rnode_178to179_bb2__22_i1469_0_reg_179_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb2__23_i1470_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i1470_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__23_i1470_0_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i1470_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i1470_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__23_i1470_1_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i1470_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__23_i1470_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i1470_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i1470_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i1470_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb2__23_i1470_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb2__23_i1470_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb2__23_i1470_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb2__23_i1470_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb2__23_i1470_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb2__23_i1470),
	.data_out(rnode_178to179_bb2__23_i1470_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb2__23_i1470_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb2__23_i1470_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb2__23_i1470_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb2__23_i1470_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb2__23_i1470_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__23_i1470_stall_in = 1'b0;
assign rnode_178to179_bb2__23_i1470_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb2__23_i1470_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__23_i1470_0_NO_SHIFT_REG = rnode_178to179_bb2__23_i1470_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb2__23_i1470_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__23_i1470_1_NO_SHIFT_REG = rnode_178to179_bb2__23_i1470_0_reg_179_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__22_i921_stall_local;
wire [31:0] local_bb2__22_i921;

assign local_bb2__22_i921 = (local_bb2__21_i920 ? local_bb2_var__u25 : rnode_177to178_bb2_add320_i1273_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i921_valid_out;
wire local_bb2__22_i921_stall_in;
 reg local_bb2__22_i921_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i922_valid_out;
wire local_bb2__23_i922_stall_in;
 reg local_bb2__23_i922_consumed_0_NO_SHIFT_REG;
wire local_bb2__23_i922_inputs_ready;
wire local_bb2__23_i922_stall_local;
wire [31:0] local_bb2__23_i922;

assign local_bb2__23_i922_inputs_ready = (rnode_177to178_bb2_c0_ene6_0_valid_out_NO_SHIFT_REG & rnode_177to178_bb2_add320_i1273_0_valid_out_2_NO_SHIFT_REG & rnode_177to178_bb2_add320_i1273_0_valid_out_3_NO_SHIFT_REG & rnode_177to178_bb2_add320_i1273_0_valid_out_1_NO_SHIFT_REG & rnode_177to178_bb2_add320_i1273_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2__23_i922 = (local_bb2__21_i920 ? rnode_177to178_bb2_add320_i1273_3_NO_SHIFT_REG : local_bb2_var__u25);
assign local_bb2__22_i921_valid_out = 1'b1;
assign local_bb2__23_i922_valid_out = 1'b1;
assign rnode_177to178_bb2_c0_ene6_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add320_i1273_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add320_i1273_0_stall_in_3_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add320_i1273_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_177to178_bb2_add320_i1273_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__22_i921_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__23_i922_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__22_i921_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i922_inputs_ready & (local_bb2__22_i921_consumed_0_NO_SHIFT_REG | ~(local_bb2__22_i921_stall_in)) & local_bb2__23_i922_stall_local);
		local_bb2__23_i922_consumed_0_NO_SHIFT_REG <= (local_bb2__23_i922_inputs_ready & (local_bb2__23_i922_consumed_0_NO_SHIFT_REG | ~(local_bb2__23_i922_stall_in)) & local_bb2__23_i922_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_shr18_i1473_stall_local;
wire [31:0] local_bb2_shr18_i1473;

assign local_bb2_shr18_i1473 = (rnode_178to179_bb2__22_i1469_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2__22_i1469_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i1469_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__22_i1469_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i1469_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i1469_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__22_i1469_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i1469_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__22_i1469_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i1469_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i1469_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i1469_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2__22_i1469_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2__22_i1469_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2__22_i1469_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2__22_i1469_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2__22_i1469_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(rnode_178to179_bb2__22_i1469_1_NO_SHIFT_REG),
	.data_out(rnode_179to180_bb2__22_i1469_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2__22_i1469_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2__22_i1469_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb2__22_i1469_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2__22_i1469_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2__22_i1469_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__22_i1469_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__22_i1469_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__22_i1469_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__22_i1469_0_NO_SHIFT_REG = rnode_179to180_bb2__22_i1469_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2__22_i1469_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__22_i1469_1_NO_SHIFT_REG = rnode_179to180_bb2__22_i1469_0_reg_180_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i1471_stall_local;
wire [31:0] local_bb2_shr16_i1471;

assign local_bb2_shr16_i1471 = (rnode_178to179_bb2__23_i1470_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2__23_i1470_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__23_i1470_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__23_i1470_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__23_i1470_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__23_i1470_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i1470_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2__23_i1470_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2__23_i1470_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2__23_i1470_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2__23_i1470_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2__23_i1470_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(rnode_178to179_bb2__23_i1470_1_NO_SHIFT_REG),
	.data_out(rnode_179to180_bb2__23_i1470_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2__23_i1470_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2__23_i1470_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb2__23_i1470_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2__23_i1470_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2__23_i1470_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__23_i1470_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__23_i1470_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__23_i1470_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__23_i1470_0_NO_SHIFT_REG = rnode_179to180_bb2__23_i1470_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2__23_i1470_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__23_i1470_1_NO_SHIFT_REG = rnode_179to180_bb2__23_i1470_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2__23_i1470_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__23_i1470_2_NO_SHIFT_REG = rnode_179to180_bb2__23_i1470_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb2__22_i921_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i921_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__22_i921_0_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i921_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i921_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__22_i921_1_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i921_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__22_i921_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i921_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i921_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__22_i921_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb2__22_i921_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb2__22_i921_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb2__22_i921_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb2__22_i921_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb2__22_i921_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb2__22_i921),
	.data_out(rnode_178to179_bb2__22_i921_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb2__22_i921_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb2__22_i921_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb2__22_i921_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb2__22_i921_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb2__22_i921_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__22_i921_stall_in = 1'b0;
assign rnode_178to179_bb2__22_i921_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb2__22_i921_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__22_i921_0_NO_SHIFT_REG = rnode_178to179_bb2__22_i921_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb2__22_i921_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__22_i921_1_NO_SHIFT_REG = rnode_178to179_bb2__22_i921_0_reg_179_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_178to179_bb2__23_i922_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i922_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__23_i922_0_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i922_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i922_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__23_i922_1_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i922_0_reg_179_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_178to179_bb2__23_i922_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i922_0_valid_out_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i922_0_stall_in_0_reg_179_NO_SHIFT_REG;
 logic rnode_178to179_bb2__23_i922_0_stall_out_reg_179_NO_SHIFT_REG;

acl_data_fifo rnode_178to179_bb2__23_i922_0_reg_179_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_178to179_bb2__23_i922_0_reg_179_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_178to179_bb2__23_i922_0_stall_in_0_reg_179_NO_SHIFT_REG),
	.valid_out(rnode_178to179_bb2__23_i922_0_valid_out_0_reg_179_NO_SHIFT_REG),
	.stall_out(rnode_178to179_bb2__23_i922_0_stall_out_reg_179_NO_SHIFT_REG),
	.data_in(local_bb2__23_i922),
	.data_out(rnode_178to179_bb2__23_i922_0_reg_179_NO_SHIFT_REG)
);

defparam rnode_178to179_bb2__23_i922_0_reg_179_fifo.DEPTH = 1;
defparam rnode_178to179_bb2__23_i922_0_reg_179_fifo.DATA_WIDTH = 32;
defparam rnode_178to179_bb2__23_i922_0_reg_179_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_178to179_bb2__23_i922_0_reg_179_fifo.IMPL = "shift_reg";

assign rnode_178to179_bb2__23_i922_0_reg_179_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__23_i922_stall_in = 1'b0;
assign rnode_178to179_bb2__23_i922_0_stall_in_0_reg_179_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb2__23_i922_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__23_i922_0_NO_SHIFT_REG = rnode_178to179_bb2__23_i922_0_reg_179_NO_SHIFT_REG;
assign rnode_178to179_bb2__23_i922_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__23_i922_1_NO_SHIFT_REG = rnode_178to179_bb2__23_i922_0_reg_179_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and19_i1474_stall_local;
wire [31:0] local_bb2_and19_i1474;

assign local_bb2_and19_i1474 = (local_bb2_shr18_i1473 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and21_i1476_stall_local;
wire [31:0] local_bb2_and21_i1476;

assign local_bb2_and21_i1476 = (rnode_179to180_bb2__22_i1469_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i1503_stall_local;
wire [31:0] local_bb2_sub_i1503;

assign local_bb2_sub_i1503 = (local_bb2_shr16_i1471 - local_bb2_shr18_i1473);

// This section implements an unregistered operation.
// 
wire local_bb2_and20_i1475_stall_local;
wire [31:0] local_bb2_and20_i1475;

assign local_bb2_and20_i1475 = (rnode_179to180_bb2__23_i1470_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and35_i1481_valid_out;
wire local_bb2_and35_i1481_stall_in;
wire local_bb2_and35_i1481_inputs_ready;
wire local_bb2_and35_i1481_stall_local;
wire [31:0] local_bb2_and35_i1481;

assign local_bb2_and35_i1481_inputs_ready = rnode_179to180_bb2__23_i1470_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and35_i1481 = (rnode_179to180_bb2__23_i1470_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb2_and35_i1481_valid_out = 1'b1;
assign rnode_179to180_bb2__23_i1470_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i1482_stall_local;
wire [31:0] local_bb2_xor_i1482;

assign local_bb2_xor_i1482 = (rnode_179to180_bb2__23_i1470_2_NO_SHIFT_REG ^ rnode_179to180_bb2__22_i1469_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shr18_i925_stall_local;
wire [31:0] local_bb2_shr18_i925;

assign local_bb2_shr18_i925 = (rnode_178to179_bb2__22_i921_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2__22_i921_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i921_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__22_i921_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i921_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i921_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__22_i921_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i921_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__22_i921_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i921_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i921_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__22_i921_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2__22_i921_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2__22_i921_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2__22_i921_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2__22_i921_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2__22_i921_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(rnode_178to179_bb2__22_i921_1_NO_SHIFT_REG),
	.data_out(rnode_179to180_bb2__22_i921_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2__22_i921_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2__22_i921_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb2__22_i921_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2__22_i921_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2__22_i921_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__22_i921_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__22_i921_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__22_i921_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__22_i921_0_NO_SHIFT_REG = rnode_179to180_bb2__22_i921_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2__22_i921_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__22_i921_1_NO_SHIFT_REG = rnode_179to180_bb2__22_i921_0_reg_180_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i923_stall_local;
wire [31:0] local_bb2_shr16_i923;

assign local_bb2_shr16_i923 = (rnode_178to179_bb2__23_i922_0_NO_SHIFT_REG >> 32'h17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2__23_i922_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__23_i922_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__23_i922_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__23_i922_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2__23_i922_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2__23_i922_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2__23_i922_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2__23_i922_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2__23_i922_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2__23_i922_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2__23_i922_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(rnode_178to179_bb2__23_i922_1_NO_SHIFT_REG),
	.data_out(rnode_179to180_bb2__23_i922_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2__23_i922_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2__23_i922_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb2__23_i922_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2__23_i922_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2__23_i922_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_178to179_bb2__23_i922_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__23_i922_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__23_i922_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__23_i922_0_NO_SHIFT_REG = rnode_179to180_bb2__23_i922_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2__23_i922_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__23_i922_1_NO_SHIFT_REG = rnode_179to180_bb2__23_i922_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2__23_i922_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2__23_i922_2_NO_SHIFT_REG = rnode_179to180_bb2__23_i922_0_reg_180_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot23_i1478_stall_local;
wire local_bb2_lnot23_i1478;

assign local_bb2_lnot23_i1478 = (local_bb2_and19_i1474 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp27_i1480_stall_local;
wire local_bb2_cmp27_i1480;

assign local_bb2_cmp27_i1480 = (local_bb2_and19_i1474 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot33_not_i1487_stall_local;
wire local_bb2_lnot33_not_i1487;

assign local_bb2_lnot33_not_i1487 = (local_bb2_and21_i1476 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or64_i1500_stall_local;
wire [31:0] local_bb2_or64_i1500;

assign local_bb2_or64_i1500 = (local_bb2_and21_i1476 << 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and68_i1504_stall_local;
wire [31:0] local_bb2_and68_i1504;

assign local_bb2_and68_i1504 = (local_bb2_sub_i1503 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_i1485_stall_local;
wire local_bb2_lnot30_i1485;

assign local_bb2_lnot30_i1485 = (local_bb2_and20_i1475 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i1497_stall_local;
wire [31:0] local_bb2_or_i1497;

assign local_bb2_or_i1497 = (local_bb2_and20_i1475 << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb2_and35_i1481_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i1481_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_and35_i1481_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i1481_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_and35_i1481_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i1481_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i1481_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i1481_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb2_and35_i1481_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb2_and35_i1481_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb2_and35_i1481_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb2_and35_i1481_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb2_and35_i1481_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb2_and35_i1481),
	.data_out(rnode_180to181_bb2_and35_i1481_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb2_and35_i1481_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb2_and35_i1481_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb2_and35_i1481_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb2_and35_i1481_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb2_and35_i1481_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and35_i1481_stall_in = 1'b0;
assign rnode_180to181_bb2_and35_i1481_0_NO_SHIFT_REG = rnode_180to181_bb2_and35_i1481_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_and35_i1481_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb2_and35_i1481_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i1483_stall_local;
wire local_bb2_cmp37_i1483;

assign local_bb2_cmp37_i1483 = ($signed(local_bb2_xor_i1482) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_xor_lobit_i1556_stall_local;
wire [31:0] local_bb2_xor_lobit_i1556;

assign local_bb2_xor_lobit_i1556 = ($signed(local_bb2_xor_i1482) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and36_lobit_i1558_stall_local;
wire [31:0] local_bb2_and36_lobit_i1558;

assign local_bb2_and36_lobit_i1558 = (local_bb2_xor_i1482 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and19_i926_stall_local;
wire [31:0] local_bb2_and19_i926;

assign local_bb2_and19_i926 = (local_bb2_shr18_i925 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and21_i928_stall_local;
wire [31:0] local_bb2_and21_i928;

assign local_bb2_and21_i928 = (rnode_179to180_bb2__22_i921_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i955_stall_local;
wire [31:0] local_bb2_sub_i955;

assign local_bb2_sub_i955 = (local_bb2_shr16_i923 - local_bb2_shr18_i925);

// This section implements an unregistered operation.
// 
wire local_bb2_and20_i927_stall_local;
wire [31:0] local_bb2_and20_i927;

assign local_bb2_and20_i927 = (rnode_179to180_bb2__23_i922_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and35_i933_valid_out;
wire local_bb2_and35_i933_stall_in;
wire local_bb2_and35_i933_inputs_ready;
wire local_bb2_and35_i933_stall_local;
wire [31:0] local_bb2_and35_i933;

assign local_bb2_and35_i933_inputs_ready = rnode_179to180_bb2__23_i922_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and35_i933 = (rnode_179to180_bb2__23_i922_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb2_and35_i933_valid_out = 1'b1;
assign rnode_179to180_bb2__23_i922_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i934_stall_local;
wire [31:0] local_bb2_xor_i934;

assign local_bb2_xor_i934 = (rnode_179to180_bb2__23_i922_2_NO_SHIFT_REG ^ rnode_179to180_bb2__22_i921_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl65_i1501_stall_local;
wire [31:0] local_bb2_shl65_i1501;

assign local_bb2_shl65_i1501 = (local_bb2_or64_i1500 | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp69_i1505_stall_local;
wire local_bb2_cmp69_i1505;

assign local_bb2_cmp69_i1505 = (local_bb2_and68_i1504 > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_not_i1489_stall_local;
wire local_bb2_lnot30_not_i1489;

assign local_bb2_lnot30_not_i1489 = (local_bb2_lnot30_i1485 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i1498_stall_local;
wire [31:0] local_bb2_shl_i1498;

assign local_bb2_shl_i1498 = (local_bb2_or_i1497 | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_and35_i1481_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i1481_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and35_i1481_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i1481_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and35_i1481_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i1481_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i1481_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i1481_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_and35_i1481_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_and35_i1481_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_and35_i1481_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_and35_i1481_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_and35_i1481_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb2_and35_i1481_0_NO_SHIFT_REG),
	.data_out(rnode_181to182_bb2_and35_i1481_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_and35_i1481_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_and35_i1481_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2_and35_i1481_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_and35_i1481_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_and35_i1481_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_and35_i1481_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and35_i1481_0_NO_SHIFT_REG = rnode_181to182_bb2_and35_i1481_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and35_i1481_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and35_i1481_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot23_i930_stall_local;
wire local_bb2_lnot23_i930;

assign local_bb2_lnot23_i930 = (local_bb2_and19_i926 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp27_i932_stall_local;
wire local_bb2_cmp27_i932;

assign local_bb2_cmp27_i932 = (local_bb2_and19_i926 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot33_not_i939_stall_local;
wire local_bb2_lnot33_not_i939;

assign local_bb2_lnot33_not_i939 = (local_bb2_and21_i928 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or64_i952_stall_local;
wire [31:0] local_bb2_or64_i952;

assign local_bb2_or64_i952 = (local_bb2_and21_i928 << 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and68_i956_stall_local;
wire [31:0] local_bb2_and68_i956;

assign local_bb2_and68_i956 = (local_bb2_sub_i955 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_i937_stall_local;
wire local_bb2_lnot30_i937;

assign local_bb2_lnot30_i937 = (local_bb2_and20_i927 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i949_stall_local;
wire [31:0] local_bb2_or_i949;

assign local_bb2_or_i949 = (local_bb2_and20_i927 << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb2_and35_i933_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i933_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_and35_i933_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i933_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_and35_i933_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i933_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i933_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_and35_i933_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb2_and35_i933_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb2_and35_i933_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb2_and35_i933_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb2_and35_i933_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb2_and35_i933_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb2_and35_i933),
	.data_out(rnode_180to181_bb2_and35_i933_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb2_and35_i933_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb2_and35_i933_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb2_and35_i933_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb2_and35_i933_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb2_and35_i933_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and35_i933_stall_in = 1'b0;
assign rnode_180to181_bb2_and35_i933_0_NO_SHIFT_REG = rnode_180to181_bb2_and35_i933_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_and35_i933_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb2_and35_i933_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i935_stall_local;
wire local_bb2_cmp37_i935;

assign local_bb2_cmp37_i935 = ($signed(local_bb2_xor_i934) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_xor_lobit_i1008_stall_local;
wire [31:0] local_bb2_xor_lobit_i1008;

assign local_bb2_xor_lobit_i1008 = ($signed(local_bb2_xor_i934) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and36_lobit_i1010_stall_local;
wire [31:0] local_bb2_and36_lobit_i1010;

assign local_bb2_and36_lobit_i1010 = (local_bb2_xor_i934 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i1471_valid_out_1;
wire local_bb2_shr16_i1471_stall_in_1;
 reg local_bb2_shr16_i1471_consumed_1_NO_SHIFT_REG;
wire local_bb2_lnot23_i1478_valid_out;
wire local_bb2_lnot23_i1478_stall_in;
 reg local_bb2_lnot23_i1478_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp27_i1480_valid_out;
wire local_bb2_cmp27_i1480_stall_in;
 reg local_bb2_cmp27_i1480_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i1506_valid_out;
wire local_bb2_align_0_i1506_stall_in;
 reg local_bb2_align_0_i1506_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i1506_inputs_ready;
wire local_bb2_align_0_i1506_stall_local;
wire [31:0] local_bb2_align_0_i1506;

assign local_bb2_align_0_i1506_inputs_ready = (rnode_178to179_bb2__22_i1469_0_valid_out_0_NO_SHIFT_REG & rnode_178to179_bb2__23_i1470_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_align_0_i1506 = (local_bb2_cmp69_i1505 ? 32'h1F : local_bb2_and68_i1504);
assign local_bb2_shr16_i1471_valid_out_1 = 1'b1;
assign local_bb2_lnot23_i1478_valid_out = 1'b1;
assign local_bb2_cmp27_i1480_valid_out = 1'b1;
assign local_bb2_align_0_i1506_valid_out = 1'b1;
assign rnode_178to179_bb2__22_i1469_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb2__23_i1470_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_shr16_i1471_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lnot23_i1478_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp27_i1480_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_align_0_i1506_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_shr16_i1471_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i1506_inputs_ready & (local_bb2_shr16_i1471_consumed_1_NO_SHIFT_REG | ~(local_bb2_shr16_i1471_stall_in_1)) & local_bb2_align_0_i1506_stall_local);
		local_bb2_lnot23_i1478_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1506_inputs_ready & (local_bb2_lnot23_i1478_consumed_0_NO_SHIFT_REG | ~(local_bb2_lnot23_i1478_stall_in)) & local_bb2_align_0_i1506_stall_local);
		local_bb2_cmp27_i1480_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1506_inputs_ready & (local_bb2_cmp27_i1480_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp27_i1480_stall_in)) & local_bb2_align_0_i1506_stall_local);
		local_bb2_align_0_i1506_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i1506_inputs_ready & (local_bb2_align_0_i1506_consumed_0_NO_SHIFT_REG | ~(local_bb2_align_0_i1506_stall_in)) & local_bb2_align_0_i1506_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_and35_i1481_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i1481_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_and35_i1481_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i1481_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_and35_i1481_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i1481_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i1481_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i1481_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_and35_i1481_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_and35_i1481_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_and35_i1481_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_and35_i1481_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_and35_i1481_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb2_and35_i1481_0_NO_SHIFT_REG),
	.data_out(rnode_182to183_bb2_and35_i1481_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_and35_i1481_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_and35_i1481_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb2_and35_i1481_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_and35_i1481_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_and35_i1481_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_and35_i1481_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and35_i1481_0_NO_SHIFT_REG = rnode_182to183_bb2_and35_i1481_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_and35_i1481_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and35_i1481_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shl65_i953_stall_local;
wire [31:0] local_bb2_shl65_i953;

assign local_bb2_shl65_i953 = (local_bb2_or64_i952 | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp69_i957_stall_local;
wire local_bb2_cmp69_i957;

assign local_bb2_cmp69_i957 = (local_bb2_and68_i956 > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_not_i941_stall_local;
wire local_bb2_lnot30_not_i941;

assign local_bb2_lnot30_not_i941 = (local_bb2_lnot30_i937 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i950_stall_local;
wire [31:0] local_bb2_shl_i950;

assign local_bb2_shl_i950 = (local_bb2_or_i949 | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_and35_i933_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i933_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and35_i933_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i933_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and35_i933_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i933_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i933_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and35_i933_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_and35_i933_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_and35_i933_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_and35_i933_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_and35_i933_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_and35_i933_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb2_and35_i933_0_NO_SHIFT_REG),
	.data_out(rnode_181to182_bb2_and35_i933_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_and35_i933_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_and35_i933_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2_and35_i933_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_and35_i933_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_and35_i933_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_and35_i933_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and35_i933_0_NO_SHIFT_REG = rnode_181to182_bb2_and35_i933_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and35_i933_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and35_i933_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2_shr16_i1471_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i1471_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_shr16_i1471_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i1471_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i1471_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_shr16_i1471_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i1471_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_shr16_i1471_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i1471_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i1471_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i1471_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2_shr16_i1471_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2_shr16_i1471_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2_shr16_i1471_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2_shr16_i1471_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2_shr16_i1471_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb2_shr16_i1471),
	.data_out(rnode_179to180_bb2_shr16_i1471_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2_shr16_i1471_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2_shr16_i1471_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb2_shr16_i1471_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2_shr16_i1471_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2_shr16_i1471_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr16_i1471_stall_in_1 = 1'b0;
assign rnode_179to180_bb2_shr16_i1471_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_shr16_i1471_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_shr16_i1471_0_NO_SHIFT_REG = rnode_179to180_bb2_shr16_i1471_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_shr16_i1471_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_shr16_i1471_1_NO_SHIFT_REG = rnode_179to180_bb2_shr16_i1471_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2_lnot23_i1478_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i1478_0_stall_in_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i1478_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i1478_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i1478_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i1478_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i1478_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i1478_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2_lnot23_i1478_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2_lnot23_i1478_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2_lnot23_i1478_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2_lnot23_i1478_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2_lnot23_i1478_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb2_lnot23_i1478),
	.data_out(rnode_179to180_bb2_lnot23_i1478_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2_lnot23_i1478_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2_lnot23_i1478_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb2_lnot23_i1478_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2_lnot23_i1478_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2_lnot23_i1478_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lnot23_i1478_stall_in = 1'b0;
assign rnode_179to180_bb2_lnot23_i1478_0_NO_SHIFT_REG = rnode_179to180_bb2_lnot23_i1478_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_lnot23_i1478_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_lnot23_i1478_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2_cmp27_i1480_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i1480_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2_cmp27_i1480_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2_cmp27_i1480_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2_cmp27_i1480_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2_cmp27_i1480_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2_cmp27_i1480_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb2_cmp27_i1480),
	.data_out(rnode_179to180_bb2_cmp27_i1480_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2_cmp27_i1480_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2_cmp27_i1480_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb2_cmp27_i1480_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2_cmp27_i1480_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2_cmp27_i1480_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp27_i1480_stall_in = 1'b0;
assign rnode_179to180_bb2_cmp27_i1480_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_cmp27_i1480_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_cmp27_i1480_0_NO_SHIFT_REG = rnode_179to180_bb2_cmp27_i1480_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_cmp27_i1480_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_cmp27_i1480_1_NO_SHIFT_REG = rnode_179to180_bb2_cmp27_i1480_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_cmp27_i1480_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_cmp27_i1480_2_NO_SHIFT_REG = rnode_179to180_bb2_cmp27_i1480_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2_align_0_i1506_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i1506_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i1506_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i1506_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i1506_3_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i1506_4_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i1506_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i1506_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2_align_0_i1506_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2_align_0_i1506_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2_align_0_i1506_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2_align_0_i1506_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2_align_0_i1506_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb2_align_0_i1506),
	.data_out(rnode_179to180_bb2_align_0_i1506_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2_align_0_i1506_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2_align_0_i1506_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb2_align_0_i1506_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2_align_0_i1506_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2_align_0_i1506_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_align_0_i1506_stall_in = 1'b0;
assign rnode_179to180_bb2_align_0_i1506_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i1506_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i1506_0_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i1506_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_align_0_i1506_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i1506_1_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i1506_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_align_0_i1506_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i1506_2_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i1506_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_align_0_i1506_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i1506_3_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i1506_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_align_0_i1506_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i1506_4_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i1506_0_reg_180_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i923_valid_out_1;
wire local_bb2_shr16_i923_stall_in_1;
 reg local_bb2_shr16_i923_consumed_1_NO_SHIFT_REG;
wire local_bb2_lnot23_i930_valid_out;
wire local_bb2_lnot23_i930_stall_in;
 reg local_bb2_lnot23_i930_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp27_i932_valid_out;
wire local_bb2_cmp27_i932_stall_in;
 reg local_bb2_cmp27_i932_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i958_valid_out;
wire local_bb2_align_0_i958_stall_in;
 reg local_bb2_align_0_i958_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i958_inputs_ready;
wire local_bb2_align_0_i958_stall_local;
wire [31:0] local_bb2_align_0_i958;

assign local_bb2_align_0_i958_inputs_ready = (rnode_178to179_bb2__22_i921_0_valid_out_0_NO_SHIFT_REG & rnode_178to179_bb2__23_i922_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_align_0_i958 = (local_bb2_cmp69_i957 ? 32'h1F : local_bb2_and68_i956);
assign local_bb2_shr16_i923_valid_out_1 = 1'b1;
assign local_bb2_lnot23_i930_valid_out = 1'b1;
assign local_bb2_cmp27_i932_valid_out = 1'b1;
assign local_bb2_align_0_i958_valid_out = 1'b1;
assign rnode_178to179_bb2__22_i921_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_178to179_bb2__23_i922_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_shr16_i923_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lnot23_i930_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp27_i932_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_align_0_i958_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_shr16_i923_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i958_inputs_ready & (local_bb2_shr16_i923_consumed_1_NO_SHIFT_REG | ~(local_bb2_shr16_i923_stall_in_1)) & local_bb2_align_0_i958_stall_local);
		local_bb2_lnot23_i930_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i958_inputs_ready & (local_bb2_lnot23_i930_consumed_0_NO_SHIFT_REG | ~(local_bb2_lnot23_i930_stall_in)) & local_bb2_align_0_i958_stall_local);
		local_bb2_cmp27_i932_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i958_inputs_ready & (local_bb2_cmp27_i932_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp27_i932_stall_in)) & local_bb2_align_0_i958_stall_local);
		local_bb2_align_0_i958_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i958_inputs_ready & (local_bb2_align_0_i958_consumed_0_NO_SHIFT_REG | ~(local_bb2_align_0_i958_stall_in)) & local_bb2_align_0_i958_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_and35_i933_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i933_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_and35_i933_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i933_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_and35_i933_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i933_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i933_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and35_i933_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_and35_i933_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_and35_i933_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_and35_i933_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_and35_i933_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_and35_i933_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb2_and35_i933_0_NO_SHIFT_REG),
	.data_out(rnode_182to183_bb2_and35_i933_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_and35_i933_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_and35_i933_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb2_and35_i933_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_and35_i933_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_and35_i933_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_and35_i933_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and35_i933_0_NO_SHIFT_REG = rnode_182to183_bb2_and35_i933_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_and35_i933_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and35_i933_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and17_i1472_stall_local;
wire [31:0] local_bb2_and17_i1472;

assign local_bb2_and17_i1472 = (rnode_179to180_bb2_shr16_i1471_0_NO_SHIFT_REG & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb2_shr16_i1471_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i1471_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb2_shr16_i1471_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i1471_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb2_shr16_i1471_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i1471_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i1471_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i1471_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb2_shr16_i1471_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb2_shr16_i1471_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb2_shr16_i1471_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb2_shr16_i1471_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb2_shr16_i1471_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_179to180_bb2_shr16_i1471_1_NO_SHIFT_REG),
	.data_out(rnode_180to182_bb2_shr16_i1471_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb2_shr16_i1471_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb2_shr16_i1471_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb2_shr16_i1471_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb2_shr16_i1471_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb2_shr16_i1471_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_shr16_i1471_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_shr16_i1471_0_NO_SHIFT_REG = rnode_180to182_bb2_shr16_i1471_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb2_shr16_i1471_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_shr16_i1471_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2__28_i1502_stall_local;
wire [31:0] local_bb2__28_i1502;

assign local_bb2__28_i1502 = (rnode_179to180_bb2_lnot23_i1478_0_NO_SHIFT_REG ? 32'h0 : local_bb2_shl65_i1501);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_i1488_stall_local;
wire local_bb2_brmerge_not_i1488;

assign local_bb2_brmerge_not_i1488 = (rnode_179to180_bb2_cmp27_i1480_0_NO_SHIFT_REG & local_bb2_lnot33_not_i1487);

// This section implements an unregistered operation.
// 
wire local_bb2_and93_i1514_stall_local;
wire [31:0] local_bb2_and93_i1514;

assign local_bb2_and93_i1514 = (rnode_179to180_bb2_align_0_i1506_0_NO_SHIFT_REG & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb2_and95_i1516_stall_local;
wire [31:0] local_bb2_and95_i1516;

assign local_bb2_and95_i1516 = (rnode_179to180_bb2_align_0_i1506_1_NO_SHIFT_REG & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and115_i1532_stall_local;
wire [31:0] local_bb2_and115_i1532;

assign local_bb2_and115_i1532 = (rnode_179to180_bb2_align_0_i1506_2_NO_SHIFT_REG & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_and130_i1538_stall_local;
wire [31:0] local_bb2_and130_i1538;

assign local_bb2_and130_i1538 = (rnode_179to180_bb2_align_0_i1506_3_NO_SHIFT_REG & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and149_i1543_stall_local;
wire [31:0] local_bb2_and149_i1543;

assign local_bb2_and149_i1543 = (rnode_179to180_bb2_align_0_i1506_4_NO_SHIFT_REG & 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2_shr16_i923_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i923_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_shr16_i923_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i923_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i923_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_shr16_i923_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i923_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_shr16_i923_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i923_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i923_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_shr16_i923_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2_shr16_i923_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2_shr16_i923_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2_shr16_i923_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2_shr16_i923_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2_shr16_i923_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb2_shr16_i923),
	.data_out(rnode_179to180_bb2_shr16_i923_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2_shr16_i923_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2_shr16_i923_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb2_shr16_i923_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2_shr16_i923_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2_shr16_i923_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr16_i923_stall_in_1 = 1'b0;
assign rnode_179to180_bb2_shr16_i923_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_shr16_i923_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_shr16_i923_0_NO_SHIFT_REG = rnode_179to180_bb2_shr16_i923_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_shr16_i923_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_shr16_i923_1_NO_SHIFT_REG = rnode_179to180_bb2_shr16_i923_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2_lnot23_i930_0_valid_out_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i930_0_stall_in_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i930_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i930_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i930_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i930_0_valid_out_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i930_0_stall_in_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_lnot23_i930_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2_lnot23_i930_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2_lnot23_i930_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2_lnot23_i930_0_stall_in_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2_lnot23_i930_0_valid_out_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2_lnot23_i930_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb2_lnot23_i930),
	.data_out(rnode_179to180_bb2_lnot23_i930_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2_lnot23_i930_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2_lnot23_i930_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb2_lnot23_i930_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2_lnot23_i930_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2_lnot23_i930_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lnot23_i930_stall_in = 1'b0;
assign rnode_179to180_bb2_lnot23_i930_0_NO_SHIFT_REG = rnode_179to180_bb2_lnot23_i930_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_lnot23_i930_0_stall_in_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_lnot23_i930_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2_cmp27_i932_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_cmp27_i932_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2_cmp27_i932_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2_cmp27_i932_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2_cmp27_i932_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2_cmp27_i932_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2_cmp27_i932_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb2_cmp27_i932),
	.data_out(rnode_179to180_bb2_cmp27_i932_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2_cmp27_i932_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2_cmp27_i932_0_reg_180_fifo.DATA_WIDTH = 1;
defparam rnode_179to180_bb2_cmp27_i932_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2_cmp27_i932_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2_cmp27_i932_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp27_i932_stall_in = 1'b0;
assign rnode_179to180_bb2_cmp27_i932_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_cmp27_i932_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_cmp27_i932_0_NO_SHIFT_REG = rnode_179to180_bb2_cmp27_i932_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_cmp27_i932_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_cmp27_i932_1_NO_SHIFT_REG = rnode_179to180_bb2_cmp27_i932_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_cmp27_i932_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_cmp27_i932_2_NO_SHIFT_REG = rnode_179to180_bb2_cmp27_i932_0_reg_180_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_179to180_bb2_align_0_i958_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i958_0_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i958_1_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i958_2_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i958_3_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i958_4_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_reg_180_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_179to180_bb2_align_0_i958_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_valid_out_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_stall_in_0_reg_180_NO_SHIFT_REG;
 logic rnode_179to180_bb2_align_0_i958_0_stall_out_reg_180_NO_SHIFT_REG;

acl_data_fifo rnode_179to180_bb2_align_0_i958_0_reg_180_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_179to180_bb2_align_0_i958_0_reg_180_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_179to180_bb2_align_0_i958_0_stall_in_0_reg_180_NO_SHIFT_REG),
	.valid_out(rnode_179to180_bb2_align_0_i958_0_valid_out_0_reg_180_NO_SHIFT_REG),
	.stall_out(rnode_179to180_bb2_align_0_i958_0_stall_out_reg_180_NO_SHIFT_REG),
	.data_in(local_bb2_align_0_i958),
	.data_out(rnode_179to180_bb2_align_0_i958_0_reg_180_NO_SHIFT_REG)
);

defparam rnode_179to180_bb2_align_0_i958_0_reg_180_fifo.DEPTH = 1;
defparam rnode_179to180_bb2_align_0_i958_0_reg_180_fifo.DATA_WIDTH = 32;
defparam rnode_179to180_bb2_align_0_i958_0_reg_180_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_179to180_bb2_align_0_i958_0_reg_180_fifo.IMPL = "shift_reg";

assign rnode_179to180_bb2_align_0_i958_0_reg_180_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_align_0_i958_stall_in = 1'b0;
assign rnode_179to180_bb2_align_0_i958_0_stall_in_0_reg_180_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i958_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i958_0_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i958_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_align_0_i958_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i958_1_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i958_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_align_0_i958_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i958_2_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i958_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_align_0_i958_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i958_3_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i958_0_reg_180_NO_SHIFT_REG;
assign rnode_179to180_bb2_align_0_i958_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_align_0_i958_4_NO_SHIFT_REG = rnode_179to180_bb2_align_0_i958_0_reg_180_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i1477_stall_local;
wire local_bb2_lnot_i1477;

assign local_bb2_lnot_i1477 = (local_bb2_and17_i1472 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_i1479_stall_local;
wire local_bb2_cmp25_i1479;

assign local_bb2_cmp25_i1479 = (local_bb2_and17_i1472 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_i1507_stall_local;
wire [31:0] local_bb2_and72_i1507;

assign local_bb2_and72_i1507 = (local_bb2__28_i1502 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i1510_stall_local;
wire [31:0] local_bb2_and75_i1510;

assign local_bb2_and75_i1510 = (local_bb2__28_i1502 & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb2_and78_i1512_stall_local;
wire [31:0] local_bb2_and78_i1512;

assign local_bb2_and78_i1512 = (local_bb2__28_i1502 & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i1518_stall_local;
wire [31:0] local_bb2_and90_i1518;

assign local_bb2_and90_i1518 = (local_bb2__28_i1502 & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and87_i1519_stall_local;
wire [31:0] local_bb2_and87_i1519;

assign local_bb2_and87_i1519 = (local_bb2__28_i1502 & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb2_and84_i1520_stall_local;
wire [31:0] local_bb2_and84_i1520;

assign local_bb2_and84_i1520 = (local_bb2__28_i1502 & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u136_stall_local;
wire [31:0] local_bb2_var__u136;

assign local_bb2_var__u136 = (local_bb2__28_i1502 & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_not_i1492_stall_local;
wire local_bb2_brmerge_not_not_i1492;

assign local_bb2_brmerge_not_not_i1492 = (local_bb2_brmerge_not_i1488 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr94_i1515_stall_local;
wire [31:0] local_bb2_shr94_i1515;

assign local_bb2_shr94_i1515 = (local_bb2__28_i1502 >> local_bb2_and93_i1514);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp96_i1517_stall_local;
wire local_bb2_cmp96_i1517;

assign local_bb2_cmp96_i1517 = (local_bb2_and95_i1516 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp116_i1533_stall_local;
wire local_bb2_cmp116_i1533;

assign local_bb2_cmp116_i1533 = (local_bb2_and115_i1532 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp131_not_i1540_stall_local;
wire local_bb2_cmp131_not_i1540;

assign local_bb2_cmp131_not_i1540 = (local_bb2_and130_i1538 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_Pivot20_i1545_stall_local;
wire local_bb2_Pivot20_i1545;

assign local_bb2_Pivot20_i1545 = (local_bb2_and149_i1543 < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_SwitchLeaf_i1546_stall_local;
wire local_bb2_SwitchLeaf_i1546;

assign local_bb2_SwitchLeaf_i1546 = (local_bb2_and149_i1543 == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and17_i924_stall_local;
wire [31:0] local_bb2_and17_i924;

assign local_bb2_and17_i924 = (rnode_179to180_bb2_shr16_i923_0_NO_SHIFT_REG & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb2_shr16_i923_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i923_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb2_shr16_i923_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i923_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb2_shr16_i923_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i923_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i923_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_shr16_i923_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb2_shr16_i923_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb2_shr16_i923_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb2_shr16_i923_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb2_shr16_i923_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb2_shr16_i923_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_179to180_bb2_shr16_i923_1_NO_SHIFT_REG),
	.data_out(rnode_180to182_bb2_shr16_i923_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb2_shr16_i923_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb2_shr16_i923_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb2_shr16_i923_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb2_shr16_i923_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb2_shr16_i923_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_179to180_bb2_shr16_i923_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_shr16_i923_0_NO_SHIFT_REG = rnode_180to182_bb2_shr16_i923_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb2_shr16_i923_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_shr16_i923_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2__28_i954_stall_local;
wire [31:0] local_bb2__28_i954;

assign local_bb2__28_i954 = (rnode_179to180_bb2_lnot23_i930_0_NO_SHIFT_REG ? 32'h0 : local_bb2_shl65_i953);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_i940_stall_local;
wire local_bb2_brmerge_not_i940;

assign local_bb2_brmerge_not_i940 = (rnode_179to180_bb2_cmp27_i932_0_NO_SHIFT_REG & local_bb2_lnot33_not_i939);

// This section implements an unregistered operation.
// 
wire local_bb2_and93_i966_stall_local;
wire [31:0] local_bb2_and93_i966;

assign local_bb2_and93_i966 = (rnode_179to180_bb2_align_0_i958_0_NO_SHIFT_REG & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb2_and95_i968_stall_local;
wire [31:0] local_bb2_and95_i968;

assign local_bb2_and95_i968 = (rnode_179to180_bb2_align_0_i958_1_NO_SHIFT_REG & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and115_i984_stall_local;
wire [31:0] local_bb2_and115_i984;

assign local_bb2_and115_i984 = (rnode_179to180_bb2_align_0_i958_2_NO_SHIFT_REG & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_and130_i990_stall_local;
wire [31:0] local_bb2_and130_i990;

assign local_bb2_and130_i990 = (rnode_179to180_bb2_align_0_i958_3_NO_SHIFT_REG & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and149_i995_stall_local;
wire [31:0] local_bb2_and149_i995;

assign local_bb2_and149_i995 = (rnode_179to180_bb2_align_0_i958_4_NO_SHIFT_REG & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i1499_stall_local;
wire [31:0] local_bb2__27_i1499;

assign local_bb2__27_i1499 = (local_bb2_lnot_i1477 ? 32'h0 : local_bb2_shl_i1498);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_not_i1484_stall_local;
wire local_bb2_cmp25_not_i1484;

assign local_bb2_cmp25_not_i1484 = (local_bb2_cmp25_i1479 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_not_i1490_stall_local;
wire local_bb2_or_cond_not_i1490;

assign local_bb2_or_cond_not_i1490 = (local_bb2_cmp25_i1479 & local_bb2_lnot30_not_i1489);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u137_stall_local;
wire local_bb2_var__u137;

assign local_bb2_var__u137 = (local_bb2_cmp25_i1479 | rnode_179to180_bb2_cmp27_i1480_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_tr_i1508_stall_local;
wire [7:0] local_bb2_and72_tr_i1508;

assign local_bb2_and72_tr_i1508 = local_bb2_and72_i1507[7:0];

// This section implements an unregistered operation.
// 
wire local_bb2_cmp76_i1511_stall_local;
wire local_bb2_cmp76_i1511;

assign local_bb2_cmp76_i1511 = (local_bb2_and75_i1510 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp79_i1513_stall_local;
wire local_bb2_cmp79_i1513;

assign local_bb2_cmp79_i1513 = (local_bb2_and78_i1512 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i1521_stall_local;
wire local_bb2_cmp91_i1521;

assign local_bb2_cmp91_i1521 = (local_bb2_and90_i1518 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp88_i1522_stall_local;
wire local_bb2_cmp88_i1522;

assign local_bb2_cmp88_i1522 = (local_bb2_and87_i1519 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp85_i1523_stall_local;
wire local_bb2_cmp85_i1523;

assign local_bb2_cmp85_i1523 = (local_bb2_and84_i1520 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u138_stall_local;
wire local_bb2_var__u138;

assign local_bb2_var__u138 = (local_bb2_var__u136 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_7_i1493_stall_local;
wire local_bb2_reduction_7_i1493;

assign local_bb2_reduction_7_i1493 = (local_bb2_cmp25_i1479 & local_bb2_brmerge_not_not_i1492);

// This section implements an unregistered operation.
// 
wire local_bb2_and142_i1542_stall_local;
wire [31:0] local_bb2_and142_i1542;

assign local_bb2_and142_i1542 = (local_bb2_shr94_i1515 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr150_i1544_stall_local;
wire [31:0] local_bb2_shr150_i1544;

assign local_bb2_shr150_i1544 = (local_bb2_shr94_i1515 >> local_bb2_and149_i1543);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u139_stall_local;
wire [31:0] local_bb2_var__u139;

assign local_bb2_var__u139 = (local_bb2_shr94_i1515 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and146_i1547_stall_local;
wire [31:0] local_bb2_and146_i1547;

assign local_bb2_and146_i1547 = (local_bb2_shr94_i1515 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i929_stall_local;
wire local_bb2_lnot_i929;

assign local_bb2_lnot_i929 = (local_bb2_and17_i924 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_i931_stall_local;
wire local_bb2_cmp25_i931;

assign local_bb2_cmp25_i931 = (local_bb2_and17_i924 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_i959_stall_local;
wire [31:0] local_bb2_and72_i959;

assign local_bb2_and72_i959 = (local_bb2__28_i954 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i962_stall_local;
wire [31:0] local_bb2_and75_i962;

assign local_bb2_and75_i962 = (local_bb2__28_i954 & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb2_and78_i964_stall_local;
wire [31:0] local_bb2_and78_i964;

assign local_bb2_and78_i964 = (local_bb2__28_i954 & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i970_stall_local;
wire [31:0] local_bb2_and90_i970;

assign local_bb2_and90_i970 = (local_bb2__28_i954 & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and87_i971_stall_local;
wire [31:0] local_bb2_and87_i971;

assign local_bb2_and87_i971 = (local_bb2__28_i954 & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb2_and84_i972_stall_local;
wire [31:0] local_bb2_and84_i972;

assign local_bb2_and84_i972 = (local_bb2__28_i954 & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u140_stall_local;
wire [31:0] local_bb2_var__u140;

assign local_bb2_var__u140 = (local_bb2__28_i954 & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_not_i944_stall_local;
wire local_bb2_brmerge_not_not_i944;

assign local_bb2_brmerge_not_not_i944 = (local_bb2_brmerge_not_i940 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr94_i967_stall_local;
wire [31:0] local_bb2_shr94_i967;

assign local_bb2_shr94_i967 = (local_bb2__28_i954 >> local_bb2_and93_i966);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp96_i969_stall_local;
wire local_bb2_cmp96_i969;

assign local_bb2_cmp96_i969 = (local_bb2_and95_i968 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp116_i985_stall_local;
wire local_bb2_cmp116_i985;

assign local_bb2_cmp116_i985 = (local_bb2_and115_i984 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp131_not_i992_stall_local;
wire local_bb2_cmp131_not_i992;

assign local_bb2_cmp131_not_i992 = (local_bb2_and130_i990 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_Pivot20_i997_stall_local;
wire local_bb2_Pivot20_i997;

assign local_bb2_Pivot20_i997 = (local_bb2_and149_i995 < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_SwitchLeaf_i998_stall_local;
wire local_bb2_SwitchLeaf_i998;

assign local_bb2_SwitchLeaf_i998 = (local_bb2_and149_i995 == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i1559_stall_local;
wire [31:0] local_bb2_add_i1559;

assign local_bb2_add_i1559 = (local_bb2__27_i1499 | local_bb2_and36_lobit_i1558);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_i1486_stall_local;
wire local_bb2_or_cond_i1486;

assign local_bb2_or_cond_i1486 = (local_bb2_lnot30_i1485 | local_bb2_cmp25_not_i1484);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i1491_stall_local;
wire local_bb2__24_i1491;

assign local_bb2__24_i1491 = (local_bb2_or_cond_not_i1490 | local_bb2_brmerge_not_i1488);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool74_i1509_stall_local;
wire [7:0] local_bb2_frombool74_i1509;

assign local_bb2_frombool74_i1509 = (local_bb2_and72_tr_i1508 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_v_i1529_stall_local;
wire local_bb2__31_v_i1529;

assign local_bb2__31_v_i1529 = (local_bb2_cmp96_i1517 ? local_bb2_cmp79_i1513 : local_bb2_cmp91_i1521);

// This section implements an unregistered operation.
// 
wire local_bb2__30_v_i1527_stall_local;
wire local_bb2__30_v_i1527;

assign local_bb2__30_v_i1527 = (local_bb2_cmp96_i1517 ? local_bb2_cmp76_i1511 : local_bb2_cmp88_i1522);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool109_i1525_stall_local;
wire [7:0] local_bb2_frombool109_i1525;

assign local_bb2_frombool109_i1525[7:1] = 7'h0;
assign local_bb2_frombool109_i1525[0] = local_bb2_cmp85_i1523;

// This section implements an unregistered operation.
// 
wire local_bb2_or107_i1524_stall_local;
wire [31:0] local_bb2_or107_i1524;

assign local_bb2_or107_i1524[31:1] = 31'h0;
assign local_bb2_or107_i1524[0] = local_bb2_var__u138;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u141_stall_local;
wire [31:0] local_bb2_var__u141;

assign local_bb2_var__u141 = (local_bb2_and146_i1547 | local_bb2_shr94_i1515);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i951_stall_local;
wire [31:0] local_bb2__27_i951;

assign local_bb2__27_i951 = (local_bb2_lnot_i929 ? 32'h0 : local_bb2_shl_i950);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_not_i936_stall_local;
wire local_bb2_cmp25_not_i936;

assign local_bb2_cmp25_not_i936 = (local_bb2_cmp25_i931 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_not_i942_stall_local;
wire local_bb2_or_cond_not_i942;

assign local_bb2_or_cond_not_i942 = (local_bb2_cmp25_i931 & local_bb2_lnot30_not_i941);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u142_stall_local;
wire local_bb2_var__u142;

assign local_bb2_var__u142 = (local_bb2_cmp25_i931 | rnode_179to180_bb2_cmp27_i932_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_tr_i960_stall_local;
wire [7:0] local_bb2_and72_tr_i960;

assign local_bb2_and72_tr_i960 = local_bb2_and72_i959[7:0];

// This section implements an unregistered operation.
// 
wire local_bb2_cmp76_i963_stall_local;
wire local_bb2_cmp76_i963;

assign local_bb2_cmp76_i963 = (local_bb2_and75_i962 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp79_i965_stall_local;
wire local_bb2_cmp79_i965;

assign local_bb2_cmp79_i965 = (local_bb2_and78_i964 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i973_stall_local;
wire local_bb2_cmp91_i973;

assign local_bb2_cmp91_i973 = (local_bb2_and90_i970 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp88_i974_stall_local;
wire local_bb2_cmp88_i974;

assign local_bb2_cmp88_i974 = (local_bb2_and87_i971 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp85_i975_stall_local;
wire local_bb2_cmp85_i975;

assign local_bb2_cmp85_i975 = (local_bb2_and84_i972 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u143_stall_local;
wire local_bb2_var__u143;

assign local_bb2_var__u143 = (local_bb2_var__u140 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_7_i945_stall_local;
wire local_bb2_reduction_7_i945;

assign local_bb2_reduction_7_i945 = (local_bb2_cmp25_i931 & local_bb2_brmerge_not_not_i944);

// This section implements an unregistered operation.
// 
wire local_bb2_and142_i994_stall_local;
wire [31:0] local_bb2_and142_i994;

assign local_bb2_and142_i994 = (local_bb2_shr94_i967 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr150_i996_stall_local;
wire [31:0] local_bb2_shr150_i996;

assign local_bb2_shr150_i996 = (local_bb2_shr94_i967 >> local_bb2_and149_i995);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u144_stall_local;
wire [31:0] local_bb2_var__u144;

assign local_bb2_var__u144 = (local_bb2_shr94_i967 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and146_i999_stall_local;
wire [31:0] local_bb2_and146_i999;

assign local_bb2_and146_i999 = (local_bb2_shr94_i967 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_8_i1494_stall_local;
wire local_bb2_reduction_8_i1494;

assign local_bb2_reduction_8_i1494 = (rnode_179to180_bb2_cmp27_i1480_1_NO_SHIFT_REG & local_bb2_or_cond_i1486);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i1530_stall_local;
wire [7:0] local_bb2__31_i1530;

assign local_bb2__31_i1530[7:1] = 7'h0;
assign local_bb2__31_i1530[0] = local_bb2__31_v_i1529;

// This section implements an unregistered operation.
// 
wire local_bb2__30_i1528_stall_local;
wire [7:0] local_bb2__30_i1528;

assign local_bb2__30_i1528[7:1] = 7'h0;
assign local_bb2__30_i1528[0] = local_bb2__30_v_i1527;

// This section implements an unregistered operation.
// 
wire local_bb2__29_i1526_stall_local;
wire [7:0] local_bb2__29_i1526;

assign local_bb2__29_i1526 = (local_bb2_cmp96_i1517 ? local_bb2_frombool74_i1509 : local_bb2_frombool109_i1525);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i1531_stall_local;
wire [31:0] local_bb2__32_i1531;

assign local_bb2__32_i1531 = (local_bb2_cmp96_i1517 ? 32'h0 : local_bb2_or107_i1524);

// This section implements an unregistered operation.
// 
wire local_bb2_or1596_i1548_stall_local;
wire [31:0] local_bb2_or1596_i1548;

assign local_bb2_or1596_i1548 = (local_bb2_var__u141 | local_bb2_and142_i1542);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i1011_stall_local;
wire [31:0] local_bb2_add_i1011;

assign local_bb2_add_i1011 = (local_bb2__27_i951 | local_bb2_and36_lobit_i1010);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_i938_stall_local;
wire local_bb2_or_cond_i938;

assign local_bb2_or_cond_i938 = (local_bb2_lnot30_i937 | local_bb2_cmp25_not_i936);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i943_stall_local;
wire local_bb2__24_i943;

assign local_bb2__24_i943 = (local_bb2_or_cond_not_i942 | local_bb2_brmerge_not_i940);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool74_i961_stall_local;
wire [7:0] local_bb2_frombool74_i961;

assign local_bb2_frombool74_i961 = (local_bb2_and72_tr_i960 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__31_v_i981_stall_local;
wire local_bb2__31_v_i981;

assign local_bb2__31_v_i981 = (local_bb2_cmp96_i969 ? local_bb2_cmp79_i965 : local_bb2_cmp91_i973);

// This section implements an unregistered operation.
// 
wire local_bb2__30_v_i979_stall_local;
wire local_bb2__30_v_i979;

assign local_bb2__30_v_i979 = (local_bb2_cmp96_i969 ? local_bb2_cmp76_i963 : local_bb2_cmp88_i974);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool109_i977_stall_local;
wire [7:0] local_bb2_frombool109_i977;

assign local_bb2_frombool109_i977[7:1] = 7'h0;
assign local_bb2_frombool109_i977[0] = local_bb2_cmp85_i975;

// This section implements an unregistered operation.
// 
wire local_bb2_or107_i976_stall_local;
wire [31:0] local_bb2_or107_i976;

assign local_bb2_or107_i976[31:1] = 31'h0;
assign local_bb2_or107_i976[0] = local_bb2_var__u143;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u145_stall_local;
wire [31:0] local_bb2_var__u145;

assign local_bb2_var__u145 = (local_bb2_and146_i999 | local_bb2_shr94_i967);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_9_i1495_stall_local;
wire local_bb2_reduction_9_i1495;

assign local_bb2_reduction_9_i1495 = (local_bb2_reduction_7_i1493 & local_bb2_reduction_8_i1494);

// This section implements an unregistered operation.
// 
wire local_bb2_or1237_i1534_stall_local;
wire [7:0] local_bb2_or1237_i1534;

assign local_bb2_or1237_i1534 = (local_bb2__30_i1528 | local_bb2__29_i1526);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i1536_stall_local;
wire [7:0] local_bb2__33_i1536;

assign local_bb2__33_i1536 = (local_bb2_cmp116_i1533 ? local_bb2__29_i1526 : local_bb2__31_i1530);

// This section implements an unregistered operation.
// 
wire local_bb2_or162_i1549_stall_local;
wire [31:0] local_bb2_or162_i1549;

assign local_bb2_or162_i1549 = (local_bb2_or1596_i1548 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_8_i946_stall_local;
wire local_bb2_reduction_8_i946;

assign local_bb2_reduction_8_i946 = (rnode_179to180_bb2_cmp27_i932_1_NO_SHIFT_REG & local_bb2_or_cond_i938);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i982_stall_local;
wire [7:0] local_bb2__31_i982;

assign local_bb2__31_i982[7:1] = 7'h0;
assign local_bb2__31_i982[0] = local_bb2__31_v_i981;

// This section implements an unregistered operation.
// 
wire local_bb2__30_i980_stall_local;
wire [7:0] local_bb2__30_i980;

assign local_bb2__30_i980[7:1] = 7'h0;
assign local_bb2__30_i980[0] = local_bb2__30_v_i979;

// This section implements an unregistered operation.
// 
wire local_bb2__29_i978_stall_local;
wire [7:0] local_bb2__29_i978;

assign local_bb2__29_i978 = (local_bb2_cmp96_i969 ? local_bb2_frombool74_i961 : local_bb2_frombool109_i977);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i983_stall_local;
wire [31:0] local_bb2__32_i983;

assign local_bb2__32_i983 = (local_bb2_cmp96_i969 ? 32'h0 : local_bb2_or107_i976);

// This section implements an unregistered operation.
// 
wire local_bb2_or1596_i1000_stall_local;
wire [31:0] local_bb2_or1596_i1000;

assign local_bb2_or1596_i1000 = (local_bb2_var__u145 | local_bb2_and142_i994);

// This section implements an unregistered operation.
// 
wire local_bb2__26_i1496_stall_local;
wire local_bb2__26_i1496;

assign local_bb2__26_i1496 = (local_bb2_reduction_9_i1495 ? local_bb2_cmp37_i1483 : local_bb2__24_i1491);

// This section implements an unregistered operation.
// 
wire local_bb2_or123_i1535_stall_local;
wire [31:0] local_bb2_or123_i1535;

assign local_bb2_or123_i1535[31:8] = 24'h0;
assign local_bb2_or123_i1535[7:0] = local_bb2_or1237_i1534;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u146_stall_local;
wire [7:0] local_bb2_var__u146;

assign local_bb2_var__u146 = (local_bb2__33_i1536 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__37_v_i1550_stall_local;
wire [31:0] local_bb2__37_v_i1550;

assign local_bb2__37_v_i1550 = (local_bb2_Pivot20_i1545 ? 32'h0 : local_bb2_or162_i1549);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_9_i947_stall_local;
wire local_bb2_reduction_9_i947;

assign local_bb2_reduction_9_i947 = (local_bb2_reduction_7_i945 & local_bb2_reduction_8_i946);

// This section implements an unregistered operation.
// 
wire local_bb2_or1237_i986_stall_local;
wire [7:0] local_bb2_or1237_i986;

assign local_bb2_or1237_i986 = (local_bb2__30_i980 | local_bb2__29_i978);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i988_stall_local;
wire [7:0] local_bb2__33_i988;

assign local_bb2__33_i988 = (local_bb2_cmp116_i985 ? local_bb2__29_i978 : local_bb2__31_i982);

// This section implements an unregistered operation.
// 
wire local_bb2_or162_i1001_stall_local;
wire [31:0] local_bb2_or162_i1001;

assign local_bb2_or162_i1001 = (local_bb2_or1596_i1000 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or124_i1537_stall_local;
wire [31:0] local_bb2_or124_i1537;

assign local_bb2_or124_i1537 = (local_bb2_cmp116_i1533 ? 32'h0 : local_bb2_or123_i1535);

// This section implements an unregistered operation.
// 
wire local_bb2_conv135_i1539_stall_local;
wire [31:0] local_bb2_conv135_i1539;

assign local_bb2_conv135_i1539[31:8] = 24'h0;
assign local_bb2_conv135_i1539[7:0] = local_bb2_var__u146;

// This section implements an unregistered operation.
// 
wire local_bb2__39_v_i1551_stall_local;
wire [31:0] local_bb2__39_v_i1551;

assign local_bb2__39_v_i1551 = (local_bb2_SwitchLeaf_i1546 ? local_bb2_var__u139 : local_bb2__37_v_i1550);

// This section implements an unregistered operation.
// 
wire local_bb2__26_i948_stall_local;
wire local_bb2__26_i948;

assign local_bb2__26_i948 = (local_bb2_reduction_9_i947 ? local_bb2_cmp37_i935 : local_bb2__24_i943);

// This section implements an unregistered operation.
// 
wire local_bb2_or123_i987_stall_local;
wire [31:0] local_bb2_or123_i987;

assign local_bb2_or123_i987[31:8] = 24'h0;
assign local_bb2_or123_i987[7:0] = local_bb2_or1237_i986;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u147_stall_local;
wire [7:0] local_bb2_var__u147;

assign local_bb2_var__u147 = (local_bb2__33_i988 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__37_v_i1002_stall_local;
wire [31:0] local_bb2__37_v_i1002;

assign local_bb2__37_v_i1002 = (local_bb2_Pivot20_i997 ? 32'h0 : local_bb2_or162_i1001);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i1552_stall_local;
wire [31:0] local_bb2_reduction_3_i1552;

assign local_bb2_reduction_3_i1552 = (local_bb2__32_i1531 | local_bb2_or124_i1537);

// This section implements an unregistered operation.
// 
wire local_bb2_or136_i1541_stall_local;
wire [31:0] local_bb2_or136_i1541;

assign local_bb2_or136_i1541 = (local_bb2_cmp131_not_i1540 ? local_bb2_conv135_i1539 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or124_i989_stall_local;
wire [31:0] local_bb2_or124_i989;

assign local_bb2_or124_i989 = (local_bb2_cmp116_i985 ? 32'h0 : local_bb2_or123_i987);

// This section implements an unregistered operation.
// 
wire local_bb2_conv135_i991_stall_local;
wire [31:0] local_bb2_conv135_i991;

assign local_bb2_conv135_i991[31:8] = 24'h0;
assign local_bb2_conv135_i991[7:0] = local_bb2_var__u147;

// This section implements an unregistered operation.
// 
wire local_bb2__39_v_i1003_stall_local;
wire [31:0] local_bb2__39_v_i1003;

assign local_bb2__39_v_i1003 = (local_bb2_SwitchLeaf_i998 ? local_bb2_var__u144 : local_bb2__37_v_i1002);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i1554_stall_local;
wire [31:0] local_bb2_reduction_5_i1554;

assign local_bb2_reduction_5_i1554 = (local_bb2_shr150_i1544 | local_bb2_reduction_3_i1552);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_4_i1553_stall_local;
wire [31:0] local_bb2_reduction_4_i1553;

assign local_bb2_reduction_4_i1553 = (local_bb2_or136_i1541 | local_bb2__39_v_i1551);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i1004_stall_local;
wire [31:0] local_bb2_reduction_3_i1004;

assign local_bb2_reduction_3_i1004 = (local_bb2__32_i983 | local_bb2_or124_i989);

// This section implements an unregistered operation.
// 
wire local_bb2_or136_i993_stall_local;
wire [31:0] local_bb2_or136_i993;

assign local_bb2_or136_i993 = (local_bb2_cmp131_not_i992 ? local_bb2_conv135_i991 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i1555_stall_local;
wire [31:0] local_bb2_reduction_6_i1555;

assign local_bb2_reduction_6_i1555 = (local_bb2_reduction_4_i1553 | local_bb2_reduction_5_i1554);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i1006_stall_local;
wire [31:0] local_bb2_reduction_5_i1006;

assign local_bb2_reduction_5_i1006 = (local_bb2_shr150_i996 | local_bb2_reduction_3_i1004);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_4_i1005_stall_local;
wire [31:0] local_bb2_reduction_4_i1005;

assign local_bb2_reduction_4_i1005 = (local_bb2_or136_i993 | local_bb2__39_v_i1003);

// This section implements an unregistered operation.
// 
wire local_bb2_xor188_i1557_stall_local;
wire [31:0] local_bb2_xor188_i1557;

assign local_bb2_xor188_i1557 = (local_bb2_reduction_6_i1555 ^ local_bb2_xor_lobit_i1556);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i1007_stall_local;
wire [31:0] local_bb2_reduction_6_i1007;

assign local_bb2_reduction_6_i1007 = (local_bb2_reduction_4_i1005 | local_bb2_reduction_5_i1006);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i1483_valid_out_1;
wire local_bb2_cmp37_i1483_stall_in_1;
 reg local_bb2_cmp37_i1483_consumed_1_NO_SHIFT_REG;
wire local_bb2__26_i1496_valid_out;
wire local_bb2__26_i1496_stall_in;
 reg local_bb2__26_i1496_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i1560_valid_out;
wire local_bb2_add192_i1560_stall_in;
 reg local_bb2_add192_i1560_consumed_0_NO_SHIFT_REG;
wire local_bb2_and17_i1472_valid_out_2;
wire local_bb2_and17_i1472_stall_in_2;
 reg local_bb2_and17_i1472_consumed_2_NO_SHIFT_REG;
wire local_bb2_var__u137_valid_out;
wire local_bb2_var__u137_stall_in;
 reg local_bb2_var__u137_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i1560_inputs_ready;
wire local_bb2_add192_i1560_stall_local;
wire [31:0] local_bb2_add192_i1560;

assign local_bb2_add192_i1560_inputs_ready = (rnode_179to180_bb2__22_i1469_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_cmp27_i1480_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_lnot23_i1478_0_valid_out_NO_SHIFT_REG & rnode_179to180_bb2__22_i1469_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb2__23_i1470_0_valid_out_2_NO_SHIFT_REG & rnode_179to180_bb2__23_i1470_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_cmp27_i1480_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb2_shr16_i1471_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_cmp27_i1480_0_valid_out_2_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i1506_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i1506_0_valid_out_4_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i1506_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i1506_0_valid_out_2_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i1506_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_add192_i1560 = (local_bb2_add_i1559 + local_bb2_xor188_i1557);
assign local_bb2_cmp37_i1483_valid_out_1 = 1'b1;
assign local_bb2__26_i1496_valid_out = 1'b1;
assign local_bb2_add192_i1560_valid_out = 1'b1;
assign local_bb2_and17_i1472_valid_out_2 = 1'b1;
assign local_bb2_var__u137_valid_out = 1'b1;
assign rnode_179to180_bb2__22_i1469_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_cmp27_i1480_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_lnot23_i1478_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__22_i1469_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__23_i1470_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__23_i1470_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_cmp27_i1480_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_shr16_i1471_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_cmp27_i1480_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i1506_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i1506_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i1506_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i1506_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i1506_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp37_i1483_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__26_i1496_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add192_i1560_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and17_i1472_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u137_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp37_i1483_consumed_1_NO_SHIFT_REG <= (local_bb2_add192_i1560_inputs_ready & (local_bb2_cmp37_i1483_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp37_i1483_stall_in_1)) & local_bb2_add192_i1560_stall_local);
		local_bb2__26_i1496_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1560_inputs_ready & (local_bb2__26_i1496_consumed_0_NO_SHIFT_REG | ~(local_bb2__26_i1496_stall_in)) & local_bb2_add192_i1560_stall_local);
		local_bb2_add192_i1560_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1560_inputs_ready & (local_bb2_add192_i1560_consumed_0_NO_SHIFT_REG | ~(local_bb2_add192_i1560_stall_in)) & local_bb2_add192_i1560_stall_local);
		local_bb2_and17_i1472_consumed_2_NO_SHIFT_REG <= (local_bb2_add192_i1560_inputs_ready & (local_bb2_and17_i1472_consumed_2_NO_SHIFT_REG | ~(local_bb2_and17_i1472_stall_in_2)) & local_bb2_add192_i1560_stall_local);
		local_bb2_var__u137_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1560_inputs_ready & (local_bb2_var__u137_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u137_stall_in)) & local_bb2_add192_i1560_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_xor188_i1009_stall_local;
wire [31:0] local_bb2_xor188_i1009;

assign local_bb2_xor188_i1009 = (local_bb2_reduction_6_i1007 ^ local_bb2_xor_lobit_i1008);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb2_cmp37_i1483_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_1_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_2_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i1483_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb2_cmp37_i1483_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb2_cmp37_i1483_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb2_cmp37_i1483_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb2_cmp37_i1483_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb2_cmp37_i1483_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_cmp37_i1483),
	.data_out(rnode_180to182_bb2_cmp37_i1483_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb2_cmp37_i1483_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb2_cmp37_i1483_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_180to182_bb2_cmp37_i1483_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb2_cmp37_i1483_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb2_cmp37_i1483_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp37_i1483_stall_in_1 = 1'b0;
assign rnode_180to182_bb2_cmp37_i1483_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_cmp37_i1483_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb2_cmp37_i1483_0_NO_SHIFT_REG = rnode_180to182_bb2_cmp37_i1483_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb2_cmp37_i1483_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb2_cmp37_i1483_1_NO_SHIFT_REG = rnode_180to182_bb2_cmp37_i1483_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb2_cmp37_i1483_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb2_cmp37_i1483_2_NO_SHIFT_REG = rnode_180to182_bb2_cmp37_i1483_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb2__26_i1496_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i1496_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i1496_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i1496_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i1496_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i1496_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i1496_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i1496_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb2__26_i1496_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb2__26_i1496_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb2__26_i1496_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb2__26_i1496_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb2__26_i1496_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb2__26_i1496),
	.data_out(rnode_180to181_bb2__26_i1496_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb2__26_i1496_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb2__26_i1496_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb2__26_i1496_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb2__26_i1496_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb2__26_i1496_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__26_i1496_stall_in = 1'b0;
assign rnode_180to181_bb2__26_i1496_0_NO_SHIFT_REG = rnode_180to181_bb2__26_i1496_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2__26_i1496_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb2__26_i1496_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb2_add192_i1560_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1560_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1560_1_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1560_2_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1560_3_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1560_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1560_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb2_add192_i1560_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb2_add192_i1560_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb2_add192_i1560_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb2_add192_i1560_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb2_add192_i1560_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb2_add192_i1560),
	.data_out(rnode_180to181_bb2_add192_i1560_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb2_add192_i1560_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb2_add192_i1560_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb2_add192_i1560_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb2_add192_i1560_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb2_add192_i1560_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add192_i1560_stall_in = 1'b0;
assign rnode_180to181_bb2_add192_i1560_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb2_add192_i1560_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_add192_i1560_0_NO_SHIFT_REG = rnode_180to181_bb2_add192_i1560_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_add192_i1560_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_add192_i1560_1_NO_SHIFT_REG = rnode_180to181_bb2_add192_i1560_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_add192_i1560_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_add192_i1560_2_NO_SHIFT_REG = rnode_180to181_bb2_add192_i1560_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_add192_i1560_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_add192_i1560_3_NO_SHIFT_REG = rnode_180to181_bb2_add192_i1560_0_reg_181_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb2_and17_i1472_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i1472_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb2_and17_i1472_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i1472_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb2_and17_i1472_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i1472_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i1472_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i1472_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb2_and17_i1472_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb2_and17_i1472_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb2_and17_i1472_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb2_and17_i1472_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb2_and17_i1472_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_and17_i1472),
	.data_out(rnode_180to182_bb2_and17_i1472_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb2_and17_i1472_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb2_and17_i1472_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb2_and17_i1472_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb2_and17_i1472_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb2_and17_i1472_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and17_i1472_stall_in_2 = 1'b0;
assign rnode_180to182_bb2_and17_i1472_0_NO_SHIFT_REG = rnode_180to182_bb2_and17_i1472_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb2_and17_i1472_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_and17_i1472_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb2_var__u137_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u137_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u137_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u137_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u137_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u137_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u137_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u137_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb2_var__u137_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb2_var__u137_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb2_var__u137_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb2_var__u137_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb2_var__u137_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb2_var__u137),
	.data_out(rnode_180to181_bb2_var__u137_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb2_var__u137_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb2_var__u137_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb2_var__u137_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb2_var__u137_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb2_var__u137_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u137_stall_in = 1'b0;
assign rnode_180to181_bb2_var__u137_0_NO_SHIFT_REG = rnode_180to181_bb2_var__u137_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_var__u137_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb2_var__u137_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i935_valid_out_1;
wire local_bb2_cmp37_i935_stall_in_1;
 reg local_bb2_cmp37_i935_consumed_1_NO_SHIFT_REG;
wire local_bb2__26_i948_valid_out;
wire local_bb2__26_i948_stall_in;
 reg local_bb2__26_i948_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i1012_valid_out;
wire local_bb2_add192_i1012_stall_in;
 reg local_bb2_add192_i1012_consumed_0_NO_SHIFT_REG;
wire local_bb2_and17_i924_valid_out_2;
wire local_bb2_and17_i924_stall_in_2;
 reg local_bb2_and17_i924_consumed_2_NO_SHIFT_REG;
wire local_bb2_var__u142_valid_out;
wire local_bb2_var__u142_stall_in;
 reg local_bb2_var__u142_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i1012_inputs_ready;
wire local_bb2_add192_i1012_stall_local;
wire [31:0] local_bb2_add192_i1012;

assign local_bb2_add192_i1012_inputs_ready = (rnode_179to180_bb2__22_i921_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_cmp27_i932_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_lnot23_i930_0_valid_out_NO_SHIFT_REG & rnode_179to180_bb2__22_i921_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb2__23_i922_0_valid_out_2_NO_SHIFT_REG & rnode_179to180_bb2__23_i922_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_cmp27_i932_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb2_shr16_i923_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_cmp27_i932_0_valid_out_2_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i958_0_valid_out_0_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i958_0_valid_out_4_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i958_0_valid_out_1_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i958_0_valid_out_2_NO_SHIFT_REG & rnode_179to180_bb2_align_0_i958_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_add192_i1012 = (local_bb2_add_i1011 + local_bb2_xor188_i1009);
assign local_bb2_cmp37_i935_valid_out_1 = 1'b1;
assign local_bb2__26_i948_valid_out = 1'b1;
assign local_bb2_add192_i1012_valid_out = 1'b1;
assign local_bb2_and17_i924_valid_out_2 = 1'b1;
assign local_bb2_var__u142_valid_out = 1'b1;
assign rnode_179to180_bb2__22_i921_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_cmp27_i932_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_lnot23_i930_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__22_i921_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__23_i922_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2__23_i922_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_cmp27_i932_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_shr16_i923_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_cmp27_i932_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i958_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i958_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i958_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i958_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_179to180_bb2_align_0_i958_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp37_i935_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__26_i948_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add192_i1012_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and17_i924_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u142_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp37_i935_consumed_1_NO_SHIFT_REG <= (local_bb2_add192_i1012_inputs_ready & (local_bb2_cmp37_i935_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp37_i935_stall_in_1)) & local_bb2_add192_i1012_stall_local);
		local_bb2__26_i948_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1012_inputs_ready & (local_bb2__26_i948_consumed_0_NO_SHIFT_REG | ~(local_bb2__26_i948_stall_in)) & local_bb2_add192_i1012_stall_local);
		local_bb2_add192_i1012_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1012_inputs_ready & (local_bb2_add192_i1012_consumed_0_NO_SHIFT_REG | ~(local_bb2_add192_i1012_stall_in)) & local_bb2_add192_i1012_stall_local);
		local_bb2_and17_i924_consumed_2_NO_SHIFT_REG <= (local_bb2_add192_i1012_inputs_ready & (local_bb2_and17_i924_consumed_2_NO_SHIFT_REG | ~(local_bb2_and17_i924_stall_in_2)) & local_bb2_add192_i1012_stall_local);
		local_bb2_var__u142_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i1012_inputs_ready & (local_bb2_var__u142_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u142_stall_in)) & local_bb2_add192_i1012_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_not_cmp37_i1589_stall_local;
wire local_bb2_not_cmp37_i1589;

assign local_bb2_not_cmp37_i1589 = (rnode_180to182_bb2_cmp37_i1483_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2__26_i1496_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i1496_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i1496_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i1496_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i1496_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i1496_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i1496_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i1496_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2__26_i1496_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2__26_i1496_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2__26_i1496_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2__26_i1496_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2__26_i1496_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb2__26_i1496_0_NO_SHIFT_REG),
	.data_out(rnode_181to182_bb2__26_i1496_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2__26_i1496_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2__26_i1496_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb2__26_i1496_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2__26_i1496_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2__26_i1496_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2__26_i1496_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__26_i1496_0_NO_SHIFT_REG = rnode_181to182_bb2__26_i1496_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2__26_i1496_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__26_i1496_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and193_i1561_valid_out;
wire local_bb2_and193_i1561_stall_in;
wire local_bb2_and193_i1561_inputs_ready;
wire local_bb2_and193_i1561_stall_local;
wire [31:0] local_bb2_and193_i1561;

assign local_bb2_and193_i1561_inputs_ready = rnode_180to181_bb2_add192_i1560_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_and193_i1561 = (rnode_180to181_bb2_add192_i1560_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb2_and193_i1561_valid_out = 1'b1;
assign rnode_180to181_bb2_add192_i1560_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and195_i1562_valid_out;
wire local_bb2_and195_i1562_stall_in;
wire local_bb2_and195_i1562_inputs_ready;
wire local_bb2_and195_i1562_stall_local;
wire [31:0] local_bb2_and195_i1562;

assign local_bb2_and195_i1562_inputs_ready = rnode_180to181_bb2_add192_i1560_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and195_i1562 = (rnode_180to181_bb2_add192_i1560_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb2_and195_i1562_valid_out = 1'b1;
assign rnode_180to181_bb2_add192_i1560_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and198_i1563_valid_out;
wire local_bb2_and198_i1563_stall_in;
wire local_bb2_and198_i1563_inputs_ready;
wire local_bb2_and198_i1563_stall_local;
wire [31:0] local_bb2_and198_i1563;

assign local_bb2_and198_i1563_inputs_ready = rnode_180to181_bb2_add192_i1560_0_valid_out_2_NO_SHIFT_REG;
assign local_bb2_and198_i1563 = (rnode_180to181_bb2_add192_i1560_2_NO_SHIFT_REG & 32'h1);
assign local_bb2_and198_i1563_valid_out = 1'b1;
assign rnode_180to181_bb2_add192_i1560_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and201_i1564_stall_local;
wire [31:0] local_bb2_and201_i1564;

assign local_bb2_and201_i1564 = (rnode_180to181_bb2_add192_i1560_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_var__u137_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u137_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u137_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u137_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u137_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u137_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u137_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u137_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_var__u137_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_var__u137_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_var__u137_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_var__u137_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_var__u137_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb2_var__u137_0_NO_SHIFT_REG),
	.data_out(rnode_181to182_bb2_var__u137_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_var__u137_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_var__u137_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb2_var__u137_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_var__u137_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_var__u137_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_var__u137_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_var__u137_0_NO_SHIFT_REG = rnode_181to182_bb2_var__u137_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_var__u137_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_var__u137_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb2_cmp37_i935_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_1_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_2_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_cmp37_i935_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb2_cmp37_i935_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb2_cmp37_i935_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb2_cmp37_i935_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb2_cmp37_i935_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb2_cmp37_i935_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_cmp37_i935),
	.data_out(rnode_180to182_bb2_cmp37_i935_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb2_cmp37_i935_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb2_cmp37_i935_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_180to182_bb2_cmp37_i935_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb2_cmp37_i935_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb2_cmp37_i935_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp37_i935_stall_in_1 = 1'b0;
assign rnode_180to182_bb2_cmp37_i935_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_cmp37_i935_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb2_cmp37_i935_0_NO_SHIFT_REG = rnode_180to182_bb2_cmp37_i935_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb2_cmp37_i935_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb2_cmp37_i935_1_NO_SHIFT_REG = rnode_180to182_bb2_cmp37_i935_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb2_cmp37_i935_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to182_bb2_cmp37_i935_2_NO_SHIFT_REG = rnode_180to182_bb2_cmp37_i935_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb2__26_i948_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i948_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i948_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i948_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i948_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i948_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i948_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2__26_i948_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb2__26_i948_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb2__26_i948_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb2__26_i948_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb2__26_i948_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb2__26_i948_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb2__26_i948),
	.data_out(rnode_180to181_bb2__26_i948_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb2__26_i948_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb2__26_i948_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb2__26_i948_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb2__26_i948_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb2__26_i948_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__26_i948_stall_in = 1'b0;
assign rnode_180to181_bb2__26_i948_0_NO_SHIFT_REG = rnode_180to181_bb2__26_i948_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2__26_i948_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb2__26_i948_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb2_add192_i1012_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1012_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1012_1_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1012_2_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1012_3_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to181_bb2_add192_i1012_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_valid_out_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_stall_in_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_add192_i1012_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb2_add192_i1012_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb2_add192_i1012_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb2_add192_i1012_0_stall_in_0_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb2_add192_i1012_0_valid_out_0_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb2_add192_i1012_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb2_add192_i1012),
	.data_out(rnode_180to181_bb2_add192_i1012_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb2_add192_i1012_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb2_add192_i1012_0_reg_181_fifo.DATA_WIDTH = 32;
defparam rnode_180to181_bb2_add192_i1012_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb2_add192_i1012_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb2_add192_i1012_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add192_i1012_stall_in = 1'b0;
assign rnode_180to181_bb2_add192_i1012_0_stall_in_0_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb2_add192_i1012_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_add192_i1012_0_NO_SHIFT_REG = rnode_180to181_bb2_add192_i1012_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_add192_i1012_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_add192_i1012_1_NO_SHIFT_REG = rnode_180to181_bb2_add192_i1012_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_add192_i1012_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_add192_i1012_2_NO_SHIFT_REG = rnode_180to181_bb2_add192_i1012_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_add192_i1012_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_add192_i1012_3_NO_SHIFT_REG = rnode_180to181_bb2_add192_i1012_0_reg_181_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_180to182_bb2_and17_i924_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i924_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb2_and17_i924_0_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i924_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_180to182_bb2_and17_i924_0_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i924_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i924_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_180to182_bb2_and17_i924_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_180to182_bb2_and17_i924_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to182_bb2_and17_i924_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to182_bb2_and17_i924_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_180to182_bb2_and17_i924_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_180to182_bb2_and17_i924_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_and17_i924),
	.data_out(rnode_180to182_bb2_and17_i924_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_180to182_bb2_and17_i924_0_reg_182_fifo.DEPTH = 2;
defparam rnode_180to182_bb2_and17_i924_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_180to182_bb2_and17_i924_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to182_bb2_and17_i924_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_180to182_bb2_and17_i924_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and17_i924_stall_in_2 = 1'b0;
assign rnode_180to182_bb2_and17_i924_0_NO_SHIFT_REG = rnode_180to182_bb2_and17_i924_0_reg_182_NO_SHIFT_REG;
assign rnode_180to182_bb2_and17_i924_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_and17_i924_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_180to181_bb2_var__u142_0_valid_out_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u142_0_stall_in_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u142_0_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u142_0_reg_181_inputs_ready_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u142_0_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u142_0_valid_out_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u142_0_stall_in_reg_181_NO_SHIFT_REG;
 logic rnode_180to181_bb2_var__u142_0_stall_out_reg_181_NO_SHIFT_REG;

acl_data_fifo rnode_180to181_bb2_var__u142_0_reg_181_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_180to181_bb2_var__u142_0_reg_181_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_180to181_bb2_var__u142_0_stall_in_reg_181_NO_SHIFT_REG),
	.valid_out(rnode_180to181_bb2_var__u142_0_valid_out_reg_181_NO_SHIFT_REG),
	.stall_out(rnode_180to181_bb2_var__u142_0_stall_out_reg_181_NO_SHIFT_REG),
	.data_in(local_bb2_var__u142),
	.data_out(rnode_180to181_bb2_var__u142_0_reg_181_NO_SHIFT_REG)
);

defparam rnode_180to181_bb2_var__u142_0_reg_181_fifo.DEPTH = 1;
defparam rnode_180to181_bb2_var__u142_0_reg_181_fifo.DATA_WIDTH = 1;
defparam rnode_180to181_bb2_var__u142_0_reg_181_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_180to181_bb2_var__u142_0_reg_181_fifo.IMPL = "shift_reg";

assign rnode_180to181_bb2_var__u142_0_reg_181_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u142_stall_in = 1'b0;
assign rnode_180to181_bb2_var__u142_0_NO_SHIFT_REG = rnode_180to181_bb2_var__u142_0_reg_181_NO_SHIFT_REG;
assign rnode_180to181_bb2_var__u142_0_stall_in_reg_181_NO_SHIFT_REG = 1'b0;
assign rnode_180to181_bb2_var__u142_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2__26_i1496_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_2_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i1496_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2__26_i1496_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2__26_i1496_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2__26_i1496_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2__26_i1496_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2__26_i1496_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb2__26_i1496_0_NO_SHIFT_REG),
	.data_out(rnode_182to183_bb2__26_i1496_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2__26_i1496_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2__26_i1496_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2__26_i1496_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2__26_i1496_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2__26_i1496_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2__26_i1496_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i1496_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i1496_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2__26_i1496_0_NO_SHIFT_REG = rnode_182to183_bb2__26_i1496_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2__26_i1496_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2__26_i1496_1_NO_SHIFT_REG = rnode_182to183_bb2__26_i1496_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2__26_i1496_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2__26_i1496_2_NO_SHIFT_REG = rnode_182to183_bb2__26_i1496_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_and193_i1561_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and193_i1561_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and193_i1561_1_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and193_i1561_2_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and193_i1561_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1561_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_and193_i1561_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_and193_i1561_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_and193_i1561_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_and193_i1561_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_and193_i1561_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_and193_i1561),
	.data_out(rnode_181to182_bb2_and193_i1561_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_and193_i1561_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_and193_i1561_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2_and193_i1561_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_and193_i1561_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_and193_i1561_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and193_i1561_stall_in = 1'b0;
assign rnode_181to182_bb2_and193_i1561_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and193_i1561_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_and193_i1561_0_NO_SHIFT_REG = rnode_181to182_bb2_and193_i1561_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and193_i1561_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_and193_i1561_1_NO_SHIFT_REG = rnode_181to182_bb2_and193_i1561_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and193_i1561_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_and193_i1561_2_NO_SHIFT_REG = rnode_181to182_bb2_and193_i1561_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_and195_i1562_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1562_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and195_i1562_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1562_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and195_i1562_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1562_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1562_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1562_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_and195_i1562_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_and195_i1562_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_and195_i1562_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_and195_i1562_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_and195_i1562_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_and195_i1562),
	.data_out(rnode_181to182_bb2_and195_i1562_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_and195_i1562_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_and195_i1562_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2_and195_i1562_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_and195_i1562_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_and195_i1562_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and195_i1562_stall_in = 1'b0;
assign rnode_181to182_bb2_and195_i1562_0_NO_SHIFT_REG = rnode_181to182_bb2_and195_i1562_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and195_i1562_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and195_i1562_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_and198_i1563_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1563_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and198_i1563_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1563_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and198_i1563_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1563_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1563_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1563_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_and198_i1563_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_and198_i1563_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_and198_i1563_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_and198_i1563_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_and198_i1563_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_and198_i1563),
	.data_out(rnode_181to182_bb2_and198_i1563_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_and198_i1563_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_and198_i1563_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2_and198_i1563_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_and198_i1563_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_and198_i1563_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and198_i1563_stall_in = 1'b0;
assign rnode_181to182_bb2_and198_i1563_0_NO_SHIFT_REG = rnode_181to182_bb2_and198_i1563_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and198_i1563_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and198_i1563_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i1565_stall_local;
wire [31:0] local_bb2_shr_i_i1565;

assign local_bb2_shr_i_i1565 = (local_bb2_and201_i1564 >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_var__u137_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u137_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u137_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u137_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u137_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u137_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u137_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u137_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_var__u137_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_var__u137_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_var__u137_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_var__u137_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_var__u137_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb2_var__u137_0_NO_SHIFT_REG),
	.data_out(rnode_182to183_bb2_var__u137_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_var__u137_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_var__u137_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_var__u137_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_var__u137_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_var__u137_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_var__u137_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_var__u137_0_NO_SHIFT_REG = rnode_182to183_bb2_var__u137_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_var__u137_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_var__u137_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_not_cmp37_i1041_stall_local;
wire local_bb2_not_cmp37_i1041;

assign local_bb2_not_cmp37_i1041 = (rnode_180to182_bb2_cmp37_i935_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2__26_i948_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i948_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i948_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i948_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i948_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i948_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i948_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__26_i948_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2__26_i948_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2__26_i948_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2__26_i948_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2__26_i948_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2__26_i948_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb2__26_i948_0_NO_SHIFT_REG),
	.data_out(rnode_181to182_bb2__26_i948_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2__26_i948_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2__26_i948_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb2__26_i948_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2__26_i948_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2__26_i948_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2__26_i948_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__26_i948_0_NO_SHIFT_REG = rnode_181to182_bb2__26_i948_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2__26_i948_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__26_i948_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and193_i1013_valid_out;
wire local_bb2_and193_i1013_stall_in;
wire local_bb2_and193_i1013_inputs_ready;
wire local_bb2_and193_i1013_stall_local;
wire [31:0] local_bb2_and193_i1013;

assign local_bb2_and193_i1013_inputs_ready = rnode_180to181_bb2_add192_i1012_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_and193_i1013 = (rnode_180to181_bb2_add192_i1012_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb2_and193_i1013_valid_out = 1'b1;
assign rnode_180to181_bb2_add192_i1012_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and195_i1014_valid_out;
wire local_bb2_and195_i1014_stall_in;
wire local_bb2_and195_i1014_inputs_ready;
wire local_bb2_and195_i1014_stall_local;
wire [31:0] local_bb2_and195_i1014;

assign local_bb2_and195_i1014_inputs_ready = rnode_180to181_bb2_add192_i1012_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and195_i1014 = (rnode_180to181_bb2_add192_i1012_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb2_and195_i1014_valid_out = 1'b1;
assign rnode_180to181_bb2_add192_i1012_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and198_i1015_valid_out;
wire local_bb2_and198_i1015_stall_in;
wire local_bb2_and198_i1015_inputs_ready;
wire local_bb2_and198_i1015_stall_local;
wire [31:0] local_bb2_and198_i1015;

assign local_bb2_and198_i1015_inputs_ready = rnode_180to181_bb2_add192_i1012_0_valid_out_2_NO_SHIFT_REG;
assign local_bb2_and198_i1015 = (rnode_180to181_bb2_add192_i1012_2_NO_SHIFT_REG & 32'h1);
assign local_bb2_and198_i1015_valid_out = 1'b1;
assign rnode_180to181_bb2_add192_i1012_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and201_i1016_stall_local;
wire [31:0] local_bb2_and201_i1016;

assign local_bb2_and201_i1016 = (rnode_180to181_bb2_add192_i1012_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_var__u142_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u142_0_stall_in_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u142_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u142_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u142_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u142_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u142_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_var__u142_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_var__u142_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_var__u142_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_var__u142_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_var__u142_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_var__u142_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(rnode_180to181_bb2_var__u142_0_NO_SHIFT_REG),
	.data_out(rnode_181to182_bb2_var__u142_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_var__u142_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_var__u142_0_reg_182_fifo.DATA_WIDTH = 1;
defparam rnode_181to182_bb2_var__u142_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_var__u142_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_var__u142_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_180to181_bb2_var__u142_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_var__u142_0_NO_SHIFT_REG = rnode_181to182_bb2_var__u142_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_var__u142_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_var__u142_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cond292_i1623_stall_local;
wire [31:0] local_bb2_cond292_i1623;

assign local_bb2_cond292_i1623 = (rnode_182to183_bb2__26_i1496_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u148_stall_local;
wire [31:0] local_bb2_var__u148;

assign local_bb2_var__u148[31:1] = 31'h0;
assign local_bb2_var__u148[0] = rnode_182to183_bb2__26_i1496_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr216_i1586_stall_local;
wire [31:0] local_bb2_shr216_i1586;

assign local_bb2_shr216_i1586 = (rnode_181to182_bb2_and193_i1561_1_NO_SHIFT_REG >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__pre_i1584_stall_local;
wire [31:0] local_bb2__pre_i1584;

assign local_bb2__pre_i1584 = (rnode_181to182_bb2_and195_i1562_0_NO_SHIFT_REG & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i1566_stall_local;
wire [31:0] local_bb2_or_i_i1566;

assign local_bb2_or_i_i1566 = (local_bb2_shr_i_i1565 | local_bb2_and201_i1564);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2__26_i948_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_2_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__26_i948_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2__26_i948_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2__26_i948_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2__26_i948_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2__26_i948_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2__26_i948_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb2__26_i948_0_NO_SHIFT_REG),
	.data_out(rnode_182to183_bb2__26_i948_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2__26_i948_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2__26_i948_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2__26_i948_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2__26_i948_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2__26_i948_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2__26_i948_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i948_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i948_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2__26_i948_0_NO_SHIFT_REG = rnode_182to183_bb2__26_i948_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2__26_i948_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2__26_i948_1_NO_SHIFT_REG = rnode_182to183_bb2__26_i948_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2__26_i948_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2__26_i948_2_NO_SHIFT_REG = rnode_182to183_bb2__26_i948_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_and193_i1013_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and193_i1013_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and193_i1013_1_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and193_i1013_2_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and193_i1013_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and193_i1013_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_and193_i1013_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_and193_i1013_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_and193_i1013_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_and193_i1013_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_and193_i1013_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_and193_i1013),
	.data_out(rnode_181to182_bb2_and193_i1013_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_and193_i1013_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_and193_i1013_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2_and193_i1013_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_and193_i1013_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_and193_i1013_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and193_i1013_stall_in = 1'b0;
assign rnode_181to182_bb2_and193_i1013_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and193_i1013_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_and193_i1013_0_NO_SHIFT_REG = rnode_181to182_bb2_and193_i1013_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and193_i1013_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_and193_i1013_1_NO_SHIFT_REG = rnode_181to182_bb2_and193_i1013_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and193_i1013_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_and193_i1013_2_NO_SHIFT_REG = rnode_181to182_bb2_and193_i1013_0_reg_182_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_and195_i1014_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1014_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and195_i1014_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1014_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and195_i1014_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1014_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1014_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and195_i1014_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_and195_i1014_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_and195_i1014_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_and195_i1014_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_and195_i1014_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_and195_i1014_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_and195_i1014),
	.data_out(rnode_181to182_bb2_and195_i1014_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_and195_i1014_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_and195_i1014_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2_and195_i1014_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_and195_i1014_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_and195_i1014_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and195_i1014_stall_in = 1'b0;
assign rnode_181to182_bb2_and195_i1014_0_NO_SHIFT_REG = rnode_181to182_bb2_and195_i1014_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and195_i1014_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and195_i1014_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2_and198_i1015_0_valid_out_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1015_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and198_i1015_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1015_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2_and198_i1015_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1015_0_valid_out_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1015_0_stall_in_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2_and198_i1015_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2_and198_i1015_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2_and198_i1015_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2_and198_i1015_0_stall_in_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2_and198_i1015_0_valid_out_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2_and198_i1015_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2_and198_i1015),
	.data_out(rnode_181to182_bb2_and198_i1015_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2_and198_i1015_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2_and198_i1015_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2_and198_i1015_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2_and198_i1015_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2_and198_i1015_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and198_i1015_stall_in = 1'b0;
assign rnode_181to182_bb2_and198_i1015_0_NO_SHIFT_REG = rnode_181to182_bb2_and198_i1015_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2_and198_i1015_0_stall_in_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and198_i1015_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i1017_stall_local;
wire [31:0] local_bb2_shr_i_i1017;

assign local_bb2_shr_i_i1017 = (local_bb2_and201_i1016 >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_var__u142_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u142_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u142_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u142_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u142_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u142_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u142_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_var__u142_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_var__u142_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_var__u142_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_var__u142_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_var__u142_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_var__u142_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(rnode_181to182_bb2_var__u142_0_NO_SHIFT_REG),
	.data_out(rnode_182to183_bb2_var__u142_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_var__u142_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_var__u142_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_var__u142_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_var__u142_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_var__u142_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2_var__u142_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_var__u142_0_NO_SHIFT_REG = rnode_182to183_bb2_var__u142_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_var__u142_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_var__u142_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext_i1633_stall_local;
wire [31:0] local_bb2_lnot_ext_i1633;

assign local_bb2_lnot_ext_i1633 = (local_bb2_var__u148 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or219_i1587_stall_local;
wire [31:0] local_bb2_or219_i1587;

assign local_bb2_or219_i1587 = (local_bb2_shr216_i1586 | rnode_181to182_bb2_and198_i1563_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool213_i1585_stall_local;
wire local_bb2_tobool213_i1585;

assign local_bb2_tobool213_i1585 = (local_bb2__pre_i1584 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shr1_i_i1567_stall_local;
wire [31:0] local_bb2_shr1_i_i1567;

assign local_bb2_shr1_i_i1567 = (local_bb2_or_i_i1566 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_cond292_i1075_stall_local;
wire [31:0] local_bb2_cond292_i1075;

assign local_bb2_cond292_i1075 = (rnode_182to183_bb2__26_i948_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u149_stall_local;
wire [31:0] local_bb2_var__u149;

assign local_bb2_var__u149[31:1] = 31'h0;
assign local_bb2_var__u149[0] = rnode_182to183_bb2__26_i948_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr216_i1038_stall_local;
wire [31:0] local_bb2_shr216_i1038;

assign local_bb2_shr216_i1038 = (rnode_181to182_bb2_and193_i1013_1_NO_SHIFT_REG >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__pre_i1036_stall_local;
wire [31:0] local_bb2__pre_i1036;

assign local_bb2__pre_i1036 = (rnode_181to182_bb2_and195_i1014_0_NO_SHIFT_REG & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i1018_stall_local;
wire [31:0] local_bb2_or_i_i1018;

assign local_bb2_or_i_i1018 = (local_bb2_shr_i_i1017 | local_bb2_and201_i1016);

// This section implements an unregistered operation.
// 
wire local_bb2__40_demorgan_i1588_stall_local;
wire local_bb2__40_demorgan_i1588;

assign local_bb2__40_demorgan_i1588 = (rnode_180to182_bb2_cmp37_i1483_0_NO_SHIFT_REG | local_bb2_tobool213_i1585);

// This section implements an unregistered operation.
// 
wire local_bb2__42_i1590_stall_local;
wire local_bb2__42_i1590;

assign local_bb2__42_i1590 = (local_bb2_tobool213_i1585 & local_bb2_not_cmp37_i1589);

// This section implements an unregistered operation.
// 
wire local_bb2_or2_i_i1568_stall_local;
wire [31:0] local_bb2_or2_i_i1568;

assign local_bb2_or2_i_i1568 = (local_bb2_shr1_i_i1567 | local_bb2_or_i_i1566);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext_i1085_stall_local;
wire [31:0] local_bb2_lnot_ext_i1085;

assign local_bb2_lnot_ext_i1085 = (local_bb2_var__u149 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or219_i1039_stall_local;
wire [31:0] local_bb2_or219_i1039;

assign local_bb2_or219_i1039 = (local_bb2_shr216_i1038 | rnode_181to182_bb2_and198_i1015_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool213_i1037_stall_local;
wire local_bb2_tobool213_i1037;

assign local_bb2_tobool213_i1037 = (local_bb2__pre_i1036 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shr1_i_i1019_stall_local;
wire [31:0] local_bb2_shr1_i_i1019;

assign local_bb2_shr1_i_i1019 = (local_bb2_or_i_i1018 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2__43_i1591_stall_local;
wire [31:0] local_bb2__43_i1591;

assign local_bb2__43_i1591 = (local_bb2__42_i1590 ? 32'h0 : local_bb2__pre_i1584);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_i1569_stall_local;
wire [31:0] local_bb2_shr3_i_i1569;

assign local_bb2_shr3_i_i1569 = (local_bb2_or2_i_i1568 >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2__40_demorgan_i1040_stall_local;
wire local_bb2__40_demorgan_i1040;

assign local_bb2__40_demorgan_i1040 = (rnode_180to182_bb2_cmp37_i935_0_NO_SHIFT_REG | local_bb2_tobool213_i1037);

// This section implements an unregistered operation.
// 
wire local_bb2__42_i1042_stall_local;
wire local_bb2__42_i1042;

assign local_bb2__42_i1042 = (local_bb2_tobool213_i1037 & local_bb2_not_cmp37_i1041);

// This section implements an unregistered operation.
// 
wire local_bb2_or2_i_i1020_stall_local;
wire [31:0] local_bb2_or2_i_i1020;

assign local_bb2_or2_i_i1020 = (local_bb2_shr1_i_i1019 | local_bb2_or_i_i1018);

// This section implements an unregistered operation.
// 
wire local_bb2_or4_i_i1570_stall_local;
wire [31:0] local_bb2_or4_i_i1570;

assign local_bb2_or4_i_i1570 = (local_bb2_shr3_i_i1569 | local_bb2_or2_i_i1568);

// This section implements an unregistered operation.
// 
wire local_bb2__43_i1043_stall_local;
wire [31:0] local_bb2__43_i1043;

assign local_bb2__43_i1043 = (local_bb2__42_i1042 ? 32'h0 : local_bb2__pre_i1036);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_i1021_stall_local;
wire [31:0] local_bb2_shr3_i_i1021;

assign local_bb2_shr3_i_i1021 = (local_bb2_or2_i_i1020 >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_shr5_i_i1571_stall_local;
wire [31:0] local_bb2_shr5_i_i1571;

assign local_bb2_shr5_i_i1571 = (local_bb2_or4_i_i1570 >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_or4_i_i1022_stall_local;
wire [31:0] local_bb2_or4_i_i1022;

assign local_bb2_or4_i_i1022 = (local_bb2_shr3_i_i1021 | local_bb2_or2_i_i1020);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_i_i1572_stall_local;
wire [31:0] local_bb2_or6_i_i1572;

assign local_bb2_or6_i_i1572 = (local_bb2_shr5_i_i1571 | local_bb2_or4_i_i1570);

// This section implements an unregistered operation.
// 
wire local_bb2_shr5_i_i1023_stall_local;
wire [31:0] local_bb2_shr5_i_i1023;

assign local_bb2_shr5_i_i1023 = (local_bb2_or4_i_i1022 >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_shr7_i_i1573_stall_local;
wire [31:0] local_bb2_shr7_i_i1573;

assign local_bb2_shr7_i_i1573 = (local_bb2_or6_i_i1572 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_masked_i_i1574_stall_local;
wire [31:0] local_bb2_or6_masked_i_i1574;

assign local_bb2_or6_masked_i_i1574 = (local_bb2_or6_i_i1572 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_i_i1024_stall_local;
wire [31:0] local_bb2_or6_i_i1024;

assign local_bb2_or6_i_i1024 = (local_bb2_shr5_i_i1023 | local_bb2_or4_i_i1022);

// This section implements an unregistered operation.
// 
wire local_bb2_neg_i_i1575_stall_local;
wire [31:0] local_bb2_neg_i_i1575;

assign local_bb2_neg_i_i1575 = (local_bb2_or6_masked_i_i1574 | local_bb2_shr7_i_i1573);

// This section implements an unregistered operation.
// 
wire local_bb2_shr7_i_i1025_stall_local;
wire [31:0] local_bb2_shr7_i_i1025;

assign local_bb2_shr7_i_i1025 = (local_bb2_or6_i_i1024 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_masked_i_i1026_stall_local;
wire [31:0] local_bb2_or6_masked_i_i1026;

assign local_bb2_or6_masked_i_i1026 = (local_bb2_or6_i_i1024 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_i1576_stall_local;
wire [31:0] local_bb2_and_i_i1576;

assign local_bb2_and_i_i1576 = (local_bb2_neg_i_i1575 ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_neg_i_i1027_stall_local;
wire [31:0] local_bb2_neg_i_i1027;

assign local_bb2_neg_i_i1027 = (local_bb2_or6_masked_i_i1026 | local_bb2_shr7_i_i1025);

// This section implements an unregistered operation.
// 
wire local_bb2__and_i_i1576_valid_out;
wire local_bb2__and_i_i1576_stall_in;
wire local_bb2__and_i_i1576_inputs_ready;
wire local_bb2__and_i_i1576_stall_local;
wire [31:0] local_bb2__and_i_i1576;

thirtysix_six_comp local_bb2__and_i_i1576_popcnt_instance (
	.data(local_bb2_and_i_i1576),
	.sum(local_bb2__and_i_i1576)
);


assign local_bb2__and_i_i1576_inputs_ready = rnode_180to181_bb2_add192_i1560_0_valid_out_3_NO_SHIFT_REG;
assign local_bb2__and_i_i1576_valid_out = 1'b1;
assign rnode_180to181_bb2_add192_i1560_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_i1028_stall_local;
wire [31:0] local_bb2_and_i_i1028;

assign local_bb2_and_i_i1028 = (local_bb2_neg_i_i1027 ^ 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2__and_i_i1576_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2__and_i_i1576_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2__and_i_i1576_1_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2__and_i_i1576_2_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2__and_i_i1576_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1576_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2__and_i_i1576_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2__and_i_i1576_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2__and_i_i1576_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2__and_i_i1576_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2__and_i_i1576_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2__and_i_i1576),
	.data_out(rnode_181to182_bb2__and_i_i1576_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2__and_i_i1576_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2__and_i_i1576_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2__and_i_i1576_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2__and_i_i1576_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2__and_i_i1576_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__and_i_i1576_stall_in = 1'b0;
assign rnode_181to182_bb2__and_i_i1576_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__and_i_i1576_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2__and_i_i1576_0_NO_SHIFT_REG = rnode_181to182_bb2__and_i_i1576_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2__and_i_i1576_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2__and_i_i1576_1_NO_SHIFT_REG = rnode_181to182_bb2__and_i_i1576_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2__and_i_i1576_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2__and_i_i1576_2_NO_SHIFT_REG = rnode_181to182_bb2__and_i_i1576_0_reg_182_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__and_i_i1028_valid_out;
wire local_bb2__and_i_i1028_stall_in;
wire local_bb2__and_i_i1028_inputs_ready;
wire local_bb2__and_i_i1028_stall_local;
wire [31:0] local_bb2__and_i_i1028;

thirtysix_six_comp local_bb2__and_i_i1028_popcnt_instance (
	.data(local_bb2_and_i_i1028),
	.sum(local_bb2__and_i_i1028)
);


assign local_bb2__and_i_i1028_inputs_ready = rnode_180to181_bb2_add192_i1012_0_valid_out_3_NO_SHIFT_REG;
assign local_bb2__and_i_i1028_valid_out = 1'b1;
assign rnode_180to181_bb2_add192_i1012_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and9_i_i1577_stall_local;
wire [31:0] local_bb2_and9_i_i1577;

assign local_bb2_and9_i_i1577 = (rnode_181to182_bb2__and_i_i1576_0_NO_SHIFT_REG & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and203_i1578_stall_local;
wire [31:0] local_bb2_and203_i1578;

assign local_bb2_and203_i1578 = (rnode_181to182_bb2__and_i_i1576_1_NO_SHIFT_REG & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_and206_i1580_stall_local;
wire [31:0] local_bb2_and206_i1580;

assign local_bb2_and206_i1580 = (rnode_181to182_bb2__and_i_i1576_2_NO_SHIFT_REG & 32'h7);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_181to182_bb2__and_i_i1028_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2__and_i_i1028_0_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2__and_i_i1028_1_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2__and_i_i1028_2_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_reg_182_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_181to182_bb2__and_i_i1028_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_valid_out_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_stall_in_0_reg_182_NO_SHIFT_REG;
 logic rnode_181to182_bb2__and_i_i1028_0_stall_out_reg_182_NO_SHIFT_REG;

acl_data_fifo rnode_181to182_bb2__and_i_i1028_0_reg_182_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_181to182_bb2__and_i_i1028_0_reg_182_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_181to182_bb2__and_i_i1028_0_stall_in_0_reg_182_NO_SHIFT_REG),
	.valid_out(rnode_181to182_bb2__and_i_i1028_0_valid_out_0_reg_182_NO_SHIFT_REG),
	.stall_out(rnode_181to182_bb2__and_i_i1028_0_stall_out_reg_182_NO_SHIFT_REG),
	.data_in(local_bb2__and_i_i1028),
	.data_out(rnode_181to182_bb2__and_i_i1028_0_reg_182_NO_SHIFT_REG)
);

defparam rnode_181to182_bb2__and_i_i1028_0_reg_182_fifo.DEPTH = 1;
defparam rnode_181to182_bb2__and_i_i1028_0_reg_182_fifo.DATA_WIDTH = 32;
defparam rnode_181to182_bb2__and_i_i1028_0_reg_182_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_181to182_bb2__and_i_i1028_0_reg_182_fifo.IMPL = "shift_reg";

assign rnode_181to182_bb2__and_i_i1028_0_reg_182_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__and_i_i1028_stall_in = 1'b0;
assign rnode_181to182_bb2__and_i_i1028_0_stall_in_0_reg_182_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__and_i_i1028_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2__and_i_i1028_0_NO_SHIFT_REG = rnode_181to182_bb2__and_i_i1028_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2__and_i_i1028_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2__and_i_i1028_1_NO_SHIFT_REG = rnode_181to182_bb2__and_i_i1028_0_reg_182_NO_SHIFT_REG;
assign rnode_181to182_bb2__and_i_i1028_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_181to182_bb2__and_i_i1028_2_NO_SHIFT_REG = rnode_181to182_bb2__and_i_i1028_0_reg_182_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_sub239_i1599_stall_local;
wire [31:0] local_bb2_sub239_i1599;

assign local_bb2_sub239_i1599 = (32'h0 - local_bb2_and9_i_i1577);

// This section implements an unregistered operation.
// 
wire local_bb2_shl204_i1579_stall_local;
wire [31:0] local_bb2_shl204_i1579;

assign local_bb2_shl204_i1579 = (rnode_181to182_bb2_and193_i1561_0_NO_SHIFT_REG << local_bb2_and203_i1578);

// This section implements an unregistered operation.
// 
wire local_bb2_and9_i_i1029_stall_local;
wire [31:0] local_bb2_and9_i_i1029;

assign local_bb2_and9_i_i1029 = (rnode_181to182_bb2__and_i_i1028_0_NO_SHIFT_REG & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and203_i1030_stall_local;
wire [31:0] local_bb2_and203_i1030;

assign local_bb2_and203_i1030 = (rnode_181to182_bb2__and_i_i1028_1_NO_SHIFT_REG & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_and206_i1032_stall_local;
wire [31:0] local_bb2_and206_i1032;

assign local_bb2_and206_i1032 = (rnode_181to182_bb2__and_i_i1028_2_NO_SHIFT_REG & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_cond244_i1600_stall_local;
wire [31:0] local_bb2_cond244_i1600;

assign local_bb2_cond244_i1600 = (rnode_180to182_bb2_cmp37_i1483_2_NO_SHIFT_REG ? local_bb2_sub239_i1599 : local_bb2__43_i1591);

// This section implements an unregistered operation.
// 
wire local_bb2_and205_i1581_stall_local;
wire [31:0] local_bb2_and205_i1581;

assign local_bb2_and205_i1581 = (local_bb2_shl204_i1579 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub239_i1051_stall_local;
wire [31:0] local_bb2_sub239_i1051;

assign local_bb2_sub239_i1051 = (32'h0 - local_bb2_and9_i_i1029);

// This section implements an unregistered operation.
// 
wire local_bb2_shl204_i1031_stall_local;
wire [31:0] local_bb2_shl204_i1031;

assign local_bb2_shl204_i1031 = (rnode_181to182_bb2_and193_i1013_0_NO_SHIFT_REG << local_bb2_and203_i1030);

// This section implements an unregistered operation.
// 
wire local_bb2_add245_i1601_stall_local;
wire [31:0] local_bb2_add245_i1601;

assign local_bb2_add245_i1601 = (local_bb2_cond244_i1600 + rnode_180to182_bb2_and17_i1472_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_fold_i1603_stall_local;
wire [31:0] local_bb2_fold_i1603;

assign local_bb2_fold_i1603 = (local_bb2_cond244_i1600 + rnode_180to182_bb2_shr16_i1471_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl207_i1582_stall_local;
wire [31:0] local_bb2_shl207_i1582;

assign local_bb2_shl207_i1582 = (local_bb2_and205_i1581 << local_bb2_and206_i1580);

// This section implements an unregistered operation.
// 
wire local_bb2_cond244_i1052_stall_local;
wire [31:0] local_bb2_cond244_i1052;

assign local_bb2_cond244_i1052 = (rnode_180to182_bb2_cmp37_i935_2_NO_SHIFT_REG ? local_bb2_sub239_i1051 : local_bb2__43_i1043);

// This section implements an unregistered operation.
// 
wire local_bb2_and205_i1033_stall_local;
wire [31:0] local_bb2_and205_i1033;

assign local_bb2_and205_i1033 = (local_bb2_shl204_i1031 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and247_i1602_stall_local;
wire [31:0] local_bb2_and247_i1602;

assign local_bb2_and247_i1602 = (local_bb2_add245_i1601 & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb2_and250_i1604_stall_local;
wire [31:0] local_bb2_and250_i1604;

assign local_bb2_and250_i1604 = (local_bb2_fold_i1603 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i1615_stall_local;
wire [31:0] local_bb2_and269_i1615;

assign local_bb2_and269_i1615 = (local_bb2_fold_i1603 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and208_i1583_stall_local;
wire [31:0] local_bb2_and208_i1583;

assign local_bb2_and208_i1583 = (local_bb2_shl207_i1582 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_add245_i1053_stall_local;
wire [31:0] local_bb2_add245_i1053;

assign local_bb2_add245_i1053 = (local_bb2_cond244_i1052 + rnode_180to182_bb2_and17_i924_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_fold_i1055_stall_local;
wire [31:0] local_bb2_fold_i1055;

assign local_bb2_fold_i1055 = (local_bb2_cond244_i1052 + rnode_180to182_bb2_shr16_i923_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl207_i1034_stall_local;
wire [31:0] local_bb2_shl207_i1034;

assign local_bb2_shl207_i1034 = (local_bb2_and205_i1033 << local_bb2_and206_i1032);

// This section implements an unregistered operation.
// 
wire local_bb2_notlhs_i1605_stall_local;
wire local_bb2_notlhs_i1605;

assign local_bb2_notlhs_i1605 = (local_bb2_and247_i1602 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_notrhs_i1606_stall_local;
wire local_bb2_notrhs_i1606;

assign local_bb2_notrhs_i1606 = (local_bb2_and250_i1604 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__44_i1592_stall_local;
wire [31:0] local_bb2__44_i1592;

assign local_bb2__44_i1592 = (local_bb2__40_demorgan_i1588 ? local_bb2_and208_i1583 : local_bb2_or219_i1587);

// This section implements an unregistered operation.
// 
wire local_bb2_and247_i1054_stall_local;
wire [31:0] local_bb2_and247_i1054;

assign local_bb2_and247_i1054 = (local_bb2_add245_i1053 & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb2_and250_i1056_stall_local;
wire [31:0] local_bb2_and250_i1056;

assign local_bb2_and250_i1056 = (local_bb2_fold_i1055 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i1067_stall_local;
wire [31:0] local_bb2_and269_i1067;

assign local_bb2_and269_i1067 = (local_bb2_fold_i1055 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and208_i1035_stall_local;
wire [31:0] local_bb2_and208_i1035;

assign local_bb2_and208_i1035 = (local_bb2_shl207_i1034 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_not__46_i1607_stall_local;
wire local_bb2_not__46_i1607;

assign local_bb2_not__46_i1607 = (local_bb2_notrhs_i1606 | local_bb2_notlhs_i1605);

// This section implements an unregistered operation.
// 
wire local_bb2__45_i1593_stall_local;
wire [31:0] local_bb2__45_i1593;

assign local_bb2__45_i1593 = (local_bb2__42_i1590 ? rnode_181to182_bb2_and193_i1561_2_NO_SHIFT_REG : local_bb2__44_i1592);

// This section implements an unregistered operation.
// 
wire local_bb2_notlhs_i1057_stall_local;
wire local_bb2_notlhs_i1057;

assign local_bb2_notlhs_i1057 = (local_bb2_and247_i1054 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_notrhs_i1058_stall_local;
wire local_bb2_notrhs_i1058;

assign local_bb2_notrhs_i1058 = (local_bb2_and250_i1056 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__44_i1044_stall_local;
wire [31:0] local_bb2__44_i1044;

assign local_bb2__44_i1044 = (local_bb2__40_demorgan_i1040 ? local_bb2_and208_i1035 : local_bb2_or219_i1039);

// This section implements an unregistered operation.
// 
wire local_bb2_and225_i1594_stall_local;
wire [31:0] local_bb2_and225_i1594;

assign local_bb2_and225_i1594 = (local_bb2__45_i1593 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i1612_stall_local;
wire [31:0] local_bb2_and270_i1612;

assign local_bb2_and270_i1612 = (local_bb2__45_i1593 & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_shr271_i1613_stall_local;
wire [31:0] local_bb2_shr271_i1613;

assign local_bb2_shr271_i1613 = (local_bb2__45_i1593 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_not__46_i1059_stall_local;
wire local_bb2_not__46_i1059;

assign local_bb2_not__46_i1059 = (local_bb2_notrhs_i1058 | local_bb2_notlhs_i1057);

// This section implements an unregistered operation.
// 
wire local_bb2__45_i1045_stall_local;
wire [31:0] local_bb2__45_i1045;

assign local_bb2__45_i1045 = (local_bb2__42_i1042 ? rnode_181to182_bb2_and193_i1013_2_NO_SHIFT_REG : local_bb2__44_i1044);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_i1595_stall_local;
wire local_bb2_cmp226_i1595;

assign local_bb2_cmp226_i1595 = (local_bb2_and225_i1594 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp296_i1627_stall_local;
wire local_bb2_cmp296_i1627;

assign local_bb2_cmp296_i1627 = (local_bb2_and270_i1612 > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp299_i1628_stall_local;
wire local_bb2_cmp299_i1628;

assign local_bb2_cmp299_i1628 = (local_bb2_and270_i1612 == 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and225_i1046_stall_local;
wire [31:0] local_bb2_and225_i1046;

assign local_bb2_and225_i1046 = (local_bb2__45_i1045 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i1064_stall_local;
wire [31:0] local_bb2_and270_i1064;

assign local_bb2_and270_i1064 = (local_bb2__45_i1045 & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_shr271_i1065_stall_local;
wire [31:0] local_bb2_shr271_i1065;

assign local_bb2_shr271_i1065 = (local_bb2__45_i1045 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_not_i1596_stall_local;
wire local_bb2_cmp226_not_i1596;

assign local_bb2_cmp226_not_i1596 = (local_bb2_cmp226_i1595 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__47_i1608_stall_local;
wire local_bb2__47_i1608;

assign local_bb2__47_i1608 = (local_bb2_cmp226_i1595 | local_bb2_not__46_i1607);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_i1047_stall_local;
wire local_bb2_cmp226_i1047;

assign local_bb2_cmp226_i1047 = (local_bb2_and225_i1046 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp296_i1079_stall_local;
wire local_bb2_cmp296_i1079;

assign local_bb2_cmp296_i1079 = (local_bb2_and270_i1064 > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i1067_valid_out;
wire local_bb2_and269_i1067_stall_in;
 reg local_bb2_and269_i1067_consumed_0_NO_SHIFT_REG;
wire local_bb2_add245_i1053_valid_out_1;
wire local_bb2_add245_i1053_stall_in_1;
 reg local_bb2_add245_i1053_consumed_1_NO_SHIFT_REG;
wire local_bb2_not__46_i1059_valid_out;
wire local_bb2_not__46_i1059_stall_in;
 reg local_bb2_not__46_i1059_consumed_0_NO_SHIFT_REG;
wire local_bb2_not_cmp37_i1041_valid_out_1;
wire local_bb2_not_cmp37_i1041_stall_in_1;
 reg local_bb2_not_cmp37_i1041_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr271_i1065_valid_out;
wire local_bb2_shr271_i1065_stall_in;
 reg local_bb2_shr271_i1065_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp226_i1047_valid_out;
wire local_bb2_cmp226_i1047_stall_in;
 reg local_bb2_cmp226_i1047_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp296_i1079_valid_out;
wire local_bb2_cmp296_i1079_stall_in;
 reg local_bb2_cmp296_i1079_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i1080_valid_out;
wire local_bb2_cmp299_i1080_stall_in;
 reg local_bb2_cmp299_i1080_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i1080_inputs_ready;
wire local_bb2_cmp299_i1080_stall_local;
wire local_bb2_cmp299_i1080;

assign local_bb2_cmp299_i1080_inputs_ready = (rnode_180to182_bb2_shr16_i923_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb2_cmp37_i935_0_valid_out_2_NO_SHIFT_REG & rnode_180to182_bb2_and17_i924_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb2_cmp37_i935_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb2_and193_i1013_0_valid_out_2_NO_SHIFT_REG & rnode_180to182_bb2_cmp37_i935_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb2_and195_i1014_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb2_and193_i1013_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb2_and198_i1015_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb2_and193_i1013_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb2__and_i_i1028_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb2__and_i_i1028_0_valid_out_2_NO_SHIFT_REG & rnode_181to182_bb2__and_i_i1028_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_cmp299_i1080 = (local_bb2_and270_i1064 == 32'h4);
assign local_bb2_and269_i1067_valid_out = 1'b1;
assign local_bb2_add245_i1053_valid_out_1 = 1'b1;
assign local_bb2_not__46_i1059_valid_out = 1'b1;
assign local_bb2_not_cmp37_i1041_valid_out_1 = 1'b1;
assign local_bb2_shr271_i1065_valid_out = 1'b1;
assign local_bb2_cmp226_i1047_valid_out = 1'b1;
assign local_bb2_cmp296_i1079_valid_out = 1'b1;
assign local_bb2_cmp299_i1080_valid_out = 1'b1;
assign rnode_180to182_bb2_shr16_i923_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_cmp37_i935_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_and17_i924_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_cmp37_i935_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and193_i1013_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_cmp37_i935_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and195_i1014_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and193_i1013_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and198_i1015_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and193_i1013_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__and_i_i1028_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__and_i_i1028_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__and_i_i1028_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_and269_i1067_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add245_i1053_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_not__46_i1059_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_not_cmp37_i1041_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr271_i1065_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp226_i1047_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp296_i1079_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp299_i1080_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_and269_i1067_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1080_inputs_ready & (local_bb2_and269_i1067_consumed_0_NO_SHIFT_REG | ~(local_bb2_and269_i1067_stall_in)) & local_bb2_cmp299_i1080_stall_local);
		local_bb2_add245_i1053_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp299_i1080_inputs_ready & (local_bb2_add245_i1053_consumed_1_NO_SHIFT_REG | ~(local_bb2_add245_i1053_stall_in_1)) & local_bb2_cmp299_i1080_stall_local);
		local_bb2_not__46_i1059_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1080_inputs_ready & (local_bb2_not__46_i1059_consumed_0_NO_SHIFT_REG | ~(local_bb2_not__46_i1059_stall_in)) & local_bb2_cmp299_i1080_stall_local);
		local_bb2_not_cmp37_i1041_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp299_i1080_inputs_ready & (local_bb2_not_cmp37_i1041_consumed_1_NO_SHIFT_REG | ~(local_bb2_not_cmp37_i1041_stall_in_1)) & local_bb2_cmp299_i1080_stall_local);
		local_bb2_shr271_i1065_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1080_inputs_ready & (local_bb2_shr271_i1065_consumed_0_NO_SHIFT_REG | ~(local_bb2_shr271_i1065_stall_in)) & local_bb2_cmp299_i1080_stall_local);
		local_bb2_cmp226_i1047_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1080_inputs_ready & (local_bb2_cmp226_i1047_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp226_i1047_stall_in)) & local_bb2_cmp299_i1080_stall_local);
		local_bb2_cmp296_i1079_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1080_inputs_ready & (local_bb2_cmp296_i1079_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp296_i1079_stall_in)) & local_bb2_cmp299_i1080_stall_local);
		local_bb2_cmp299_i1080_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i1080_inputs_ready & (local_bb2_cmp299_i1080_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp299_i1080_stall_in)) & local_bb2_cmp299_i1080_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_and269_i1615_valid_out;
wire local_bb2_and269_i1615_stall_in;
 reg local_bb2_and269_i1615_consumed_0_NO_SHIFT_REG;
wire local_bb2_add245_i1601_valid_out_1;
wire local_bb2_add245_i1601_stall_in_1;
 reg local_bb2_add245_i1601_consumed_1_NO_SHIFT_REG;
wire local_bb2_brmerge12_i1597_valid_out;
wire local_bb2_brmerge12_i1597_stall_in;
 reg local_bb2_brmerge12_i1597_consumed_0_NO_SHIFT_REG;
wire local_bb2_shr271_i1613_valid_out;
wire local_bb2_shr271_i1613_stall_in;
 reg local_bb2_shr271_i1613_consumed_0_NO_SHIFT_REG;
wire local_bb2__47_i1608_valid_out;
wire local_bb2__47_i1608_stall_in;
 reg local_bb2__47_i1608_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp296_i1627_valid_out;
wire local_bb2_cmp296_i1627_stall_in;
 reg local_bb2_cmp296_i1627_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i1628_valid_out;
wire local_bb2_cmp299_i1628_stall_in;
 reg local_bb2_cmp299_i1628_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp226_not_i1596_valid_out_1;
wire local_bb2_cmp226_not_i1596_stall_in_1;
 reg local_bb2_cmp226_not_i1596_consumed_1_NO_SHIFT_REG;
wire local_bb2_brmerge12_i1597_inputs_ready;
wire local_bb2_brmerge12_i1597_stall_local;
wire local_bb2_brmerge12_i1597;

assign local_bb2_brmerge12_i1597_inputs_ready = (rnode_180to182_bb2_shr16_i1471_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb2_cmp37_i1483_0_valid_out_2_NO_SHIFT_REG & rnode_180to182_bb2_and17_i1472_0_valid_out_NO_SHIFT_REG & rnode_180to182_bb2_cmp37_i1483_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb2_and193_i1561_0_valid_out_2_NO_SHIFT_REG & rnode_180to182_bb2_cmp37_i1483_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb2_and195_i1562_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb2_and193_i1561_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb2_and198_i1563_0_valid_out_NO_SHIFT_REG & rnode_181to182_bb2_and193_i1561_0_valid_out_0_NO_SHIFT_REG & rnode_181to182_bb2__and_i_i1576_0_valid_out_1_NO_SHIFT_REG & rnode_181to182_bb2__and_i_i1576_0_valid_out_2_NO_SHIFT_REG & rnode_181to182_bb2__and_i_i1576_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_brmerge12_i1597 = (local_bb2_cmp226_not_i1596 | local_bb2_not_cmp37_i1589);
assign local_bb2_and269_i1615_valid_out = 1'b1;
assign local_bb2_add245_i1601_valid_out_1 = 1'b1;
assign local_bb2_brmerge12_i1597_valid_out = 1'b1;
assign local_bb2_shr271_i1613_valid_out = 1'b1;
assign local_bb2__47_i1608_valid_out = 1'b1;
assign local_bb2_cmp296_i1627_valid_out = 1'b1;
assign local_bb2_cmp299_i1628_valid_out = 1'b1;
assign local_bb2_cmp226_not_i1596_valid_out_1 = 1'b1;
assign rnode_180to182_bb2_shr16_i1471_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_cmp37_i1483_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_and17_i1472_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_cmp37_i1483_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and193_i1561_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_180to182_bb2_cmp37_i1483_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and195_i1562_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and193_i1561_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and198_i1563_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2_and193_i1561_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__and_i_i1576_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__and_i_i1576_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_181to182_bb2__and_i_i1576_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_and269_i1615_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add245_i1601_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_brmerge12_i1597_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr271_i1613_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__47_i1608_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp296_i1627_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp299_i1628_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp226_not_i1596_consumed_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_and269_i1615_consumed_0_NO_SHIFT_REG <= (local_bb2_brmerge12_i1597_inputs_ready & (local_bb2_and269_i1615_consumed_0_NO_SHIFT_REG | ~(local_bb2_and269_i1615_stall_in)) & local_bb2_brmerge12_i1597_stall_local);
		local_bb2_add245_i1601_consumed_1_NO_SHIFT_REG <= (local_bb2_brmerge12_i1597_inputs_ready & (local_bb2_add245_i1601_consumed_1_NO_SHIFT_REG | ~(local_bb2_add245_i1601_stall_in_1)) & local_bb2_brmerge12_i1597_stall_local);
		local_bb2_brmerge12_i1597_consumed_0_NO_SHIFT_REG <= (local_bb2_brmerge12_i1597_inputs_ready & (local_bb2_brmerge12_i1597_consumed_0_NO_SHIFT_REG | ~(local_bb2_brmerge12_i1597_stall_in)) & local_bb2_brmerge12_i1597_stall_local);
		local_bb2_shr271_i1613_consumed_0_NO_SHIFT_REG <= (local_bb2_brmerge12_i1597_inputs_ready & (local_bb2_shr271_i1613_consumed_0_NO_SHIFT_REG | ~(local_bb2_shr271_i1613_stall_in)) & local_bb2_brmerge12_i1597_stall_local);
		local_bb2__47_i1608_consumed_0_NO_SHIFT_REG <= (local_bb2_brmerge12_i1597_inputs_ready & (local_bb2__47_i1608_consumed_0_NO_SHIFT_REG | ~(local_bb2__47_i1608_stall_in)) & local_bb2_brmerge12_i1597_stall_local);
		local_bb2_cmp296_i1627_consumed_0_NO_SHIFT_REG <= (local_bb2_brmerge12_i1597_inputs_ready & (local_bb2_cmp296_i1627_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp296_i1627_stall_in)) & local_bb2_brmerge12_i1597_stall_local);
		local_bb2_cmp299_i1628_consumed_0_NO_SHIFT_REG <= (local_bb2_brmerge12_i1597_inputs_ready & (local_bb2_cmp299_i1628_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp299_i1628_stall_in)) & local_bb2_brmerge12_i1597_stall_local);
		local_bb2_cmp226_not_i1596_consumed_1_NO_SHIFT_REG <= (local_bb2_brmerge12_i1597_inputs_ready & (local_bb2_cmp226_not_i1596_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp226_not_i1596_stall_in_1)) & local_bb2_brmerge12_i1597_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_and269_i1067_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1067_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_and269_i1067_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1067_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_and269_i1067_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1067_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1067_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1067_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_and269_i1067_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_and269_i1067_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_and269_i1067_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_and269_i1067_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_and269_i1067_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_and269_i1067),
	.data_out(rnode_182to183_bb2_and269_i1067_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_and269_i1067_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_and269_i1067_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb2_and269_i1067_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_and269_i1067_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_and269_i1067_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and269_i1067_stall_in = 1'b0;
assign rnode_182to183_bb2_and269_i1067_0_NO_SHIFT_REG = rnode_182to183_bb2_and269_i1067_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_and269_i1067_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and269_i1067_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_add245_i1053_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1053_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_add245_i1053_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1053_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_add245_i1053_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1053_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1053_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1053_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_add245_i1053_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_add245_i1053_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_add245_i1053_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_add245_i1053_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_add245_i1053_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_add245_i1053),
	.data_out(rnode_182to183_bb2_add245_i1053_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_add245_i1053_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_add245_i1053_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb2_add245_i1053_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_add245_i1053_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_add245_i1053_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add245_i1053_stall_in_1 = 1'b0;
assign rnode_182to183_bb2_add245_i1053_0_NO_SHIFT_REG = rnode_182to183_bb2_add245_i1053_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_add245_i1053_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_add245_i1053_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_not__46_i1059_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not__46_i1059_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not__46_i1059_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not__46_i1059_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not__46_i1059_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not__46_i1059_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not__46_i1059_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not__46_i1059_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_not__46_i1059_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_not__46_i1059_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_not__46_i1059_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_not__46_i1059_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_not__46_i1059_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_not__46_i1059),
	.data_out(rnode_182to183_bb2_not__46_i1059_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_not__46_i1059_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_not__46_i1059_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_not__46_i1059_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_not__46_i1059_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_not__46_i1059_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not__46_i1059_stall_in = 1'b0;
assign rnode_182to183_bb2_not__46_i1059_0_NO_SHIFT_REG = rnode_182to183_bb2_not__46_i1059_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_not__46_i1059_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_not__46_i1059_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_not_cmp37_i1041_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not_cmp37_i1041_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not_cmp37_i1041_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not_cmp37_i1041_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not_cmp37_i1041_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_not_cmp37_i1041_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_not_cmp37_i1041_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_not_cmp37_i1041_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_not_cmp37_i1041_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_not_cmp37_i1041),
	.data_out(rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not_cmp37_i1041_stall_in_1 = 1'b0;
assign rnode_182to183_bb2_not_cmp37_i1041_0_NO_SHIFT_REG = rnode_182to183_bb2_not_cmp37_i1041_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_not_cmp37_i1041_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_not_cmp37_i1041_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_shr271_i1065_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1065_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_shr271_i1065_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1065_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_shr271_i1065_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1065_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1065_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1065_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_shr271_i1065_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_shr271_i1065_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_shr271_i1065_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_shr271_i1065_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_shr271_i1065_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_shr271_i1065),
	.data_out(rnode_182to183_bb2_shr271_i1065_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_shr271_i1065_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_shr271_i1065_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb2_shr271_i1065_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_shr271_i1065_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_shr271_i1065_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr271_i1065_stall_in = 1'b0;
assign rnode_182to183_bb2_shr271_i1065_0_NO_SHIFT_REG = rnode_182to183_bb2_shr271_i1065_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_shr271_i1065_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_shr271_i1065_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_cmp226_i1047_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_i1047_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_cmp226_i1047_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_cmp226_i1047_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_cmp226_i1047_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_cmp226_i1047_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_cmp226_i1047_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_cmp226_i1047),
	.data_out(rnode_182to183_bb2_cmp226_i1047_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_cmp226_i1047_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_cmp226_i1047_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_cmp226_i1047_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_cmp226_i1047_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_cmp226_i1047_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp226_i1047_stall_in = 1'b0;
assign rnode_182to183_bb2_cmp226_i1047_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp226_i1047_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2_cmp226_i1047_0_NO_SHIFT_REG = rnode_182to183_bb2_cmp226_i1047_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_cmp226_i1047_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2_cmp226_i1047_1_NO_SHIFT_REG = rnode_182to183_bb2_cmp226_i1047_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_cmp296_i1079_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1079_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1079_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1079_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1079_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1079_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1079_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1079_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_cmp296_i1079_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_cmp296_i1079_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_cmp296_i1079_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_cmp296_i1079_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_cmp296_i1079_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_cmp296_i1079),
	.data_out(rnode_182to183_bb2_cmp296_i1079_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_cmp296_i1079_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_cmp296_i1079_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_cmp296_i1079_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_cmp296_i1079_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_cmp296_i1079_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp296_i1079_stall_in = 1'b0;
assign rnode_182to183_bb2_cmp296_i1079_0_NO_SHIFT_REG = rnode_182to183_bb2_cmp296_i1079_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_cmp296_i1079_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp296_i1079_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_cmp299_i1080_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1080_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1080_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1080_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1080_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1080_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1080_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1080_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_cmp299_i1080_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_cmp299_i1080_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_cmp299_i1080_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_cmp299_i1080_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_cmp299_i1080_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_cmp299_i1080),
	.data_out(rnode_182to183_bb2_cmp299_i1080_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_cmp299_i1080_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_cmp299_i1080_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_cmp299_i1080_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_cmp299_i1080_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_cmp299_i1080_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp299_i1080_stall_in = 1'b0;
assign rnode_182to183_bb2_cmp299_i1080_0_NO_SHIFT_REG = rnode_182to183_bb2_cmp299_i1080_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_cmp299_i1080_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp299_i1080_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_and269_i1615_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1615_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_and269_i1615_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1615_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_and269_i1615_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1615_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1615_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_and269_i1615_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_and269_i1615_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_and269_i1615_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_and269_i1615_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_and269_i1615_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_and269_i1615_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_and269_i1615),
	.data_out(rnode_182to183_bb2_and269_i1615_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_and269_i1615_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_and269_i1615_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb2_and269_i1615_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_and269_i1615_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_and269_i1615_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and269_i1615_stall_in = 1'b0;
assign rnode_182to183_bb2_and269_i1615_0_NO_SHIFT_REG = rnode_182to183_bb2_and269_i1615_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_and269_i1615_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and269_i1615_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_add245_i1601_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1601_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_add245_i1601_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1601_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_add245_i1601_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1601_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1601_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_add245_i1601_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_add245_i1601_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_add245_i1601_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_add245_i1601_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_add245_i1601_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_add245_i1601_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_add245_i1601),
	.data_out(rnode_182to183_bb2_add245_i1601_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_add245_i1601_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_add245_i1601_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb2_add245_i1601_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_add245_i1601_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_add245_i1601_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add245_i1601_stall_in_1 = 1'b0;
assign rnode_182to183_bb2_add245_i1601_0_NO_SHIFT_REG = rnode_182to183_bb2_add245_i1601_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_add245_i1601_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_add245_i1601_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_brmerge12_i1597_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_brmerge12_i1597_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_brmerge12_i1597_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_brmerge12_i1597_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_brmerge12_i1597_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_brmerge12_i1597_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_brmerge12_i1597_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_brmerge12_i1597_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_brmerge12_i1597_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_brmerge12_i1597_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_brmerge12_i1597_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_brmerge12_i1597_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_brmerge12_i1597_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_brmerge12_i1597),
	.data_out(rnode_182to183_bb2_brmerge12_i1597_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_brmerge12_i1597_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_brmerge12_i1597_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_brmerge12_i1597_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_brmerge12_i1597_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_brmerge12_i1597_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_brmerge12_i1597_stall_in = 1'b0;
assign rnode_182to183_bb2_brmerge12_i1597_0_NO_SHIFT_REG = rnode_182to183_bb2_brmerge12_i1597_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_brmerge12_i1597_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_brmerge12_i1597_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_shr271_i1613_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1613_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_shr271_i1613_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1613_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_182to183_bb2_shr271_i1613_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1613_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1613_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_shr271_i1613_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_shr271_i1613_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_shr271_i1613_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_shr271_i1613_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_shr271_i1613_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_shr271_i1613_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_shr271_i1613),
	.data_out(rnode_182to183_bb2_shr271_i1613_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_shr271_i1613_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_shr271_i1613_0_reg_183_fifo.DATA_WIDTH = 32;
defparam rnode_182to183_bb2_shr271_i1613_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_shr271_i1613_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_shr271_i1613_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr271_i1613_stall_in = 1'b0;
assign rnode_182to183_bb2_shr271_i1613_0_NO_SHIFT_REG = rnode_182to183_bb2_shr271_i1613_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_shr271_i1613_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_shr271_i1613_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2__47_i1608_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_1_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_valid_out_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_stall_in_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2__47_i1608_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2__47_i1608_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2__47_i1608_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2__47_i1608_0_stall_in_0_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2__47_i1608_0_valid_out_0_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2__47_i1608_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2__47_i1608),
	.data_out(rnode_182to183_bb2__47_i1608_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2__47_i1608_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2__47_i1608_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2__47_i1608_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2__47_i1608_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2__47_i1608_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__47_i1608_stall_in = 1'b0;
assign rnode_182to183_bb2__47_i1608_0_stall_in_0_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__47_i1608_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2__47_i1608_0_NO_SHIFT_REG = rnode_182to183_bb2__47_i1608_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2__47_i1608_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_182to183_bb2__47_i1608_1_NO_SHIFT_REG = rnode_182to183_bb2__47_i1608_0_reg_183_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_cmp296_i1627_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1627_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1627_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1627_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1627_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1627_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1627_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp296_i1627_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_cmp296_i1627_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_cmp296_i1627_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_cmp296_i1627_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_cmp296_i1627_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_cmp296_i1627_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_cmp296_i1627),
	.data_out(rnode_182to183_bb2_cmp296_i1627_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_cmp296_i1627_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_cmp296_i1627_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_cmp296_i1627_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_cmp296_i1627_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_cmp296_i1627_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp296_i1627_stall_in = 1'b0;
assign rnode_182to183_bb2_cmp296_i1627_0_NO_SHIFT_REG = rnode_182to183_bb2_cmp296_i1627_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_cmp296_i1627_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp296_i1627_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_cmp299_i1628_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1628_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1628_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1628_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1628_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1628_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1628_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp299_i1628_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_cmp299_i1628_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_cmp299_i1628_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_cmp299_i1628_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_cmp299_i1628_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_cmp299_i1628_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_cmp299_i1628),
	.data_out(rnode_182to183_bb2_cmp299_i1628_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_cmp299_i1628_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_cmp299_i1628_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_cmp299_i1628_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_cmp299_i1628_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_cmp299_i1628_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp299_i1628_stall_in = 1'b0;
assign rnode_182to183_bb2_cmp299_i1628_0_NO_SHIFT_REG = rnode_182to183_bb2_cmp299_i1628_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_cmp299_i1628_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp299_i1628_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_182to183_bb2_cmp226_not_i1596_0_valid_out_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_not_i1596_0_stall_in_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_not_i1596_0_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_inputs_ready_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_not_i1596_0_valid_out_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_not_i1596_0_stall_in_reg_183_NO_SHIFT_REG;
 logic rnode_182to183_bb2_cmp226_not_i1596_0_stall_out_reg_183_NO_SHIFT_REG;

acl_data_fifo rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_182to183_bb2_cmp226_not_i1596_0_stall_in_reg_183_NO_SHIFT_REG),
	.valid_out(rnode_182to183_bb2_cmp226_not_i1596_0_valid_out_reg_183_NO_SHIFT_REG),
	.stall_out(rnode_182to183_bb2_cmp226_not_i1596_0_stall_out_reg_183_NO_SHIFT_REG),
	.data_in(local_bb2_cmp226_not_i1596),
	.data_out(rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_NO_SHIFT_REG)
);

defparam rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_fifo.DEPTH = 1;
defparam rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_fifo.DATA_WIDTH = 1;
defparam rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_fifo.IMPL = "shift_reg";

assign rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp226_not_i1596_stall_in_1 = 1'b0;
assign rnode_182to183_bb2_cmp226_not_i1596_0_NO_SHIFT_REG = rnode_182to183_bb2_cmp226_not_i1596_0_reg_183_NO_SHIFT_REG;
assign rnode_182to183_bb2_cmp226_not_i1596_0_stall_in_reg_183_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp226_not_i1596_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shl273_i1068_stall_local;
wire [31:0] local_bb2_shl273_i1068;

assign local_bb2_shl273_i1068 = (rnode_182to183_bb2_and269_i1067_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp258_i1061_stall_local;
wire local_bb2_cmp258_i1061;

assign local_bb2_cmp258_i1061 = ($signed(rnode_182to183_bb2_add245_i1053_0_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb2_and272_i1066_stall_local;
wire [31:0] local_bb2_and272_i1066;

assign local_bb2_and272_i1066 = (rnode_182to183_bb2_shr271_i1065_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_not_i1048_stall_local;
wire local_bb2_cmp226_not_i1048;

assign local_bb2_cmp226_not_i1048 = (rnode_182to183_bb2_cmp226_i1047_0_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__47_i1060_stall_local;
wire local_bb2__47_i1060;

assign local_bb2__47_i1060 = (rnode_182to183_bb2_cmp226_i1047_1_NO_SHIFT_REG | rnode_182to183_bb2_not__46_i1059_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp29649_i1083_stall_local;
wire [31:0] local_bb2_cmp29649_i1083;

assign local_bb2_cmp29649_i1083[31:1] = 31'h0;
assign local_bb2_cmp29649_i1083[0] = rnode_182to183_bb2_cmp296_i1079_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_conv300_i1081_stall_local;
wire [31:0] local_bb2_conv300_i1081;

assign local_bb2_conv300_i1081[31:1] = 31'h0;
assign local_bb2_conv300_i1081[0] = rnode_182to183_bb2_cmp299_i1080_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shl273_i1616_stall_local;
wire [31:0] local_bb2_shl273_i1616;

assign local_bb2_shl273_i1616 = (rnode_182to183_bb2_and269_i1615_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp258_i1609_stall_local;
wire local_bb2_cmp258_i1609;

assign local_bb2_cmp258_i1609 = ($signed(rnode_182to183_bb2_add245_i1601_0_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb2_resultSign_0_i1598_stall_local;
wire [31:0] local_bb2_resultSign_0_i1598;

assign local_bb2_resultSign_0_i1598 = (rnode_182to183_bb2_brmerge12_i1597_0_NO_SHIFT_REG ? rnode_182to183_bb2_and35_i1481_0_NO_SHIFT_REG : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_and272_i1614_stall_local;
wire [31:0] local_bb2_and272_i1614;

assign local_bb2_and272_i1614 = (rnode_182to183_bb2_shr271_i1613_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u150_valid_out;
wire local_bb2_var__u150_stall_in;
wire local_bb2_var__u150_inputs_ready;
wire local_bb2_var__u150_stall_local;
wire [31:0] local_bb2_var__u150;

assign local_bb2_var__u150_inputs_ready = rnode_182to183_bb2__47_i1608_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_var__u150[31:1] = 31'h0;
assign local_bb2_var__u150[0] = rnode_182to183_bb2__47_i1608_1_NO_SHIFT_REG;
assign local_bb2_var__u150_valid_out = 1'b1;
assign rnode_182to183_bb2__47_i1608_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp29649_i1631_stall_local;
wire [31:0] local_bb2_cmp29649_i1631;

assign local_bb2_cmp29649_i1631[31:1] = 31'h0;
assign local_bb2_cmp29649_i1631[0] = rnode_182to183_bb2_cmp296_i1627_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_conv300_i1629_stall_local;
wire [31:0] local_bb2_conv300_i1629;

assign local_bb2_conv300_i1629[31:1] = 31'h0;
assign local_bb2_conv300_i1629[0] = rnode_182to183_bb2_cmp299_i1628_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_or274_i1069_stall_local;
wire [31:0] local_bb2_or274_i1069;

assign local_bb2_or274_i1069 = (local_bb2_and272_i1066 | local_bb2_shl273_i1068);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge12_i1049_stall_local;
wire local_bb2_brmerge12_i1049;

assign local_bb2_brmerge12_i1049 = (local_bb2_cmp226_not_i1048 | rnode_182to183_bb2_not_cmp37_i1041_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot262__i1062_stall_local;
wire local_bb2_lnot262__i1062;

assign local_bb2_lnot262__i1062 = (local_bb2_cmp258_i1061 & local_bb2_cmp226_not_i1048);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u151_stall_local;
wire [31:0] local_bb2_var__u151;

assign local_bb2_var__u151[31:1] = 31'h0;
assign local_bb2_var__u151[0] = local_bb2__47_i1060;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot262__i1610_stall_local;
wire local_bb2_lnot262__i1610;

assign local_bb2_lnot262__i1610 = (local_bb2_cmp258_i1609 & rnode_182to183_bb2_cmp226_not_i1596_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_or274_i1617_stall_local;
wire [31:0] local_bb2_or274_i1617;

assign local_bb2_or274_i1617 = (local_bb2_and272_i1614 | local_bb2_shl273_i1616);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb2_var__u150_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u150_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_var__u150_0_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u150_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_var__u150_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u150_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u150_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u150_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb2_var__u150_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb2_var__u150_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb2_var__u150_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb2_var__u150_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb2_var__u150_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb2_var__u150),
	.data_out(rnode_183to184_bb2_var__u150_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb2_var__u150_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb2_var__u150_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb2_var__u150_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb2_var__u150_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb2_var__u150_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u150_stall_in = 1'b0;
assign rnode_183to184_bb2_var__u150_0_NO_SHIFT_REG = rnode_183to184_bb2_var__u150_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb2_var__u150_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_var__u150_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_resultSign_0_i1050_stall_local;
wire [31:0] local_bb2_resultSign_0_i1050;

assign local_bb2_resultSign_0_i1050 = (local_bb2_brmerge12_i1049 ? rnode_182to183_bb2_and35_i933_0_NO_SHIFT_REG : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or2662_i1063_stall_local;
wire local_bb2_or2662_i1063;

assign local_bb2_or2662_i1063 = (rnode_182to183_bb2_var__u142_0_NO_SHIFT_REG | local_bb2_lnot262__i1062);

// This section implements an unregistered operation.
// 
wire local_bb2_or2662_i1611_stall_local;
wire local_bb2_or2662_i1611;

assign local_bb2_or2662_i1611 = (rnode_182to183_bb2_var__u137_0_NO_SHIFT_REG | local_bb2_lnot262__i1610);

// This section implements an unregistered operation.
// 
wire local_bb2_or275_i1618_stall_local;
wire [31:0] local_bb2_or275_i1618;

assign local_bb2_or275_i1618 = (local_bb2_or274_i1617 | local_bb2_resultSign_0_i1598);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext314_i1635_stall_local;
wire [31:0] local_bb2_lnot_ext314_i1635;

assign local_bb2_lnot_ext314_i1635 = (rnode_183to184_bb2_var__u150_0_NO_SHIFT_REG ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or275_i1070_stall_local;
wire [31:0] local_bb2_or275_i1070;

assign local_bb2_or275_i1070 = (local_bb2_or274_i1069 | local_bb2_resultSign_0_i1050);

// This section implements an unregistered operation.
// 
wire local_bb2_or2804_i1071_stall_local;
wire local_bb2_or2804_i1071;

assign local_bb2_or2804_i1071 = (local_bb2__47_i1060 | local_bb2_or2662_i1063);

// This section implements an unregistered operation.
// 
wire local_bb2_or2875_i1073_stall_local;
wire local_bb2_or2875_i1073;

assign local_bb2_or2875_i1073 = (local_bb2_or2662_i1063 | rnode_182to183_bb2__26_i948_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u152_stall_local;
wire [31:0] local_bb2_var__u152;

assign local_bb2_var__u152[31:1] = 31'h0;
assign local_bb2_var__u152[0] = local_bb2_or2662_i1063;

// This section implements an unregistered operation.
// 
wire local_bb2_or2804_i1619_stall_local;
wire local_bb2_or2804_i1619;

assign local_bb2_or2804_i1619 = (rnode_182to183_bb2__47_i1608_0_NO_SHIFT_REG | local_bb2_or2662_i1611);

// This section implements an unregistered operation.
// 
wire local_bb2_or2875_i1621_stall_local;
wire local_bb2_or2875_i1621;

assign local_bb2_or2875_i1621 = (local_bb2_or2662_i1611 | rnode_182to183_bb2__26_i1496_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u153_stall_local;
wire [31:0] local_bb2_var__u153;

assign local_bb2_var__u153[31:1] = 31'h0;
assign local_bb2_var__u153[0] = local_bb2_or2662_i1611;

// This section implements an unregistered operation.
// 
wire local_bb2_cond282_i1072_stall_local;
wire [31:0] local_bb2_cond282_i1072;

assign local_bb2_cond282_i1072 = (local_bb2_or2804_i1071 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond289_i1074_stall_local;
wire [31:0] local_bb2_cond289_i1074;

assign local_bb2_cond289_i1074 = (local_bb2_or2875_i1073 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext310_i1086_stall_local;
wire [31:0] local_bb2_lnot_ext310_i1086;

assign local_bb2_lnot_ext310_i1086 = (local_bb2_var__u152 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cond282_i1620_stall_local;
wire [31:0] local_bb2_cond282_i1620;

assign local_bb2_cond282_i1620 = (local_bb2_or2804_i1619 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond289_i1622_stall_local;
wire [31:0] local_bb2_cond289_i1622;

assign local_bb2_cond289_i1622 = (local_bb2_or2875_i1621 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext310_i1634_stall_local;
wire [31:0] local_bb2_lnot_ext310_i1634;

assign local_bb2_lnot_ext310_i1634 = (local_bb2_var__u153 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and293_i1076_stall_local;
wire [31:0] local_bb2_and293_i1076;

assign local_bb2_and293_i1076 = (local_bb2_cond282_i1072 & local_bb2_or275_i1070);

// This section implements an unregistered operation.
// 
wire local_bb2_or294_i1077_stall_local;
wire [31:0] local_bb2_or294_i1077;

assign local_bb2_or294_i1077 = (local_bb2_cond289_i1074 | local_bb2_cond292_i1075);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i1088_stall_local;
wire [31:0] local_bb2_reduction_0_i1088;

assign local_bb2_reduction_0_i1088 = (local_bb2_lnot_ext310_i1086 & local_bb2_lnot_ext_i1085);

// This section implements an unregistered operation.
// 
wire local_bb2_and293_i1624_stall_local;
wire [31:0] local_bb2_and293_i1624;

assign local_bb2_and293_i1624 = (local_bb2_cond282_i1620 & local_bb2_or275_i1618);

// This section implements an unregistered operation.
// 
wire local_bb2_or294_i1625_stall_local;
wire [31:0] local_bb2_or294_i1625;

assign local_bb2_or294_i1625 = (local_bb2_cond289_i1622 | local_bb2_cond292_i1623);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i1636_stall_local;
wire [31:0] local_bb2_reduction_0_i1636;

assign local_bb2_reduction_0_i1636 = (local_bb2_lnot_ext310_i1634 & local_bb2_lnot_ext_i1633);

// This section implements an unregistered operation.
// 
wire local_bb2_and302_i1082_stall_local;
wire [31:0] local_bb2_and302_i1082;

assign local_bb2_and302_i1082 = (local_bb2_conv300_i1081 & local_bb2_and293_i1076);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i1078_stall_local;
wire [31:0] local_bb2_or295_i1078;

assign local_bb2_or295_i1078 = (local_bb2_or294_i1077 | local_bb2_and293_i1076);

// This section implements an unregistered operation.
// 
wire local_bb2_and302_i1630_stall_local;
wire [31:0] local_bb2_and302_i1630;

assign local_bb2_and302_i1630 = (local_bb2_conv300_i1629 & local_bb2_and293_i1624);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i1626_stall_local;
wire [31:0] local_bb2_or295_i1626;

assign local_bb2_or295_i1626 = (local_bb2_or294_i1625 | local_bb2_and293_i1624);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i1078_valid_out;
wire local_bb2_or295_i1078_stall_in;
 reg local_bb2_or295_i1078_consumed_0_NO_SHIFT_REG;
wire local_bb2_var__u151_valid_out;
wire local_bb2_var__u151_stall_in;
 reg local_bb2_var__u151_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i1084_valid_out;
wire local_bb2_lor_ext_i1084_stall_in;
 reg local_bb2_lor_ext_i1084_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i1088_valid_out;
wire local_bb2_reduction_0_i1088_stall_in;
 reg local_bb2_reduction_0_i1088_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i1084_inputs_ready;
wire local_bb2_lor_ext_i1084_stall_local;
wire [31:0] local_bb2_lor_ext_i1084;

assign local_bb2_lor_ext_i1084_inputs_ready = (rnode_182to183_bb2_and35_i933_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_not_cmp37_i1041_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_and269_i1067_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_add245_i1053_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_var__u142_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2__26_i948_0_valid_out_0_NO_SHIFT_REG & rnode_182to183_bb2__26_i948_0_valid_out_1_NO_SHIFT_REG & rnode_182to183_bb2_cmp226_i1047_0_valid_out_1_NO_SHIFT_REG & rnode_182to183_bb2_not__46_i1059_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_shr271_i1065_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2__26_i948_0_valid_out_2_NO_SHIFT_REG & rnode_182to183_bb2_cmp226_i1047_0_valid_out_0_NO_SHIFT_REG & rnode_182to183_bb2_cmp296_i1079_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_cmp299_i1080_0_valid_out_NO_SHIFT_REG);
assign local_bb2_lor_ext_i1084 = (local_bb2_cmp29649_i1083 | local_bb2_and302_i1082);
assign local_bb2_or295_i1078_valid_out = 1'b1;
assign local_bb2_var__u151_valid_out = 1'b1;
assign local_bb2_lor_ext_i1084_valid_out = 1'b1;
assign local_bb2_reduction_0_i1088_valid_out = 1'b1;
assign rnode_182to183_bb2_and35_i933_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_not_cmp37_i1041_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and269_i1067_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_add245_i1053_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_var__u142_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i948_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i948_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp226_i1047_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_not__46_i1059_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_shr271_i1065_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i948_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp226_i1047_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp296_i1079_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp299_i1080_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_or295_i1078_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u151_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_lor_ext_i1084_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i1088_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_or295_i1078_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1084_inputs_ready & (local_bb2_or295_i1078_consumed_0_NO_SHIFT_REG | ~(local_bb2_or295_i1078_stall_in)) & local_bb2_lor_ext_i1084_stall_local);
		local_bb2_var__u151_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1084_inputs_ready & (local_bb2_var__u151_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u151_stall_in)) & local_bb2_lor_ext_i1084_stall_local);
		local_bb2_lor_ext_i1084_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1084_inputs_ready & (local_bb2_lor_ext_i1084_consumed_0_NO_SHIFT_REG | ~(local_bb2_lor_ext_i1084_stall_in)) & local_bb2_lor_ext_i1084_stall_local);
		local_bb2_reduction_0_i1088_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1084_inputs_ready & (local_bb2_reduction_0_i1088_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i1088_stall_in)) & local_bb2_lor_ext_i1084_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_or295_i1626_valid_out;
wire local_bb2_or295_i1626_stall_in;
 reg local_bb2_or295_i1626_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i1632_valid_out;
wire local_bb2_lor_ext_i1632_stall_in;
 reg local_bb2_lor_ext_i1632_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i1636_valid_out;
wire local_bb2_reduction_0_i1636_stall_in;
 reg local_bb2_reduction_0_i1636_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i1632_inputs_ready;
wire local_bb2_lor_ext_i1632_stall_local;
wire [31:0] local_bb2_lor_ext_i1632;

assign local_bb2_lor_ext_i1632_inputs_ready = (rnode_182to183_bb2_brmerge12_i1597_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_and35_i1481_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_and269_i1615_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_add245_i1601_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_cmp226_not_i1596_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_var__u137_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2__47_i1608_0_valid_out_0_NO_SHIFT_REG & rnode_182to183_bb2__26_i1496_0_valid_out_0_NO_SHIFT_REG & rnode_182to183_bb2__26_i1496_0_valid_out_1_NO_SHIFT_REG & rnode_182to183_bb2_shr271_i1613_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2__26_i1496_0_valid_out_2_NO_SHIFT_REG & rnode_182to183_bb2_cmp296_i1627_0_valid_out_NO_SHIFT_REG & rnode_182to183_bb2_cmp299_i1628_0_valid_out_NO_SHIFT_REG);
assign local_bb2_lor_ext_i1632 = (local_bb2_cmp29649_i1631 | local_bb2_and302_i1630);
assign local_bb2_or295_i1626_valid_out = 1'b1;
assign local_bb2_lor_ext_i1632_valid_out = 1'b1;
assign local_bb2_reduction_0_i1636_valid_out = 1'b1;
assign rnode_182to183_bb2_brmerge12_i1597_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and35_i1481_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_and269_i1615_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_add245_i1601_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp226_not_i1596_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_var__u137_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__47_i1608_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i1496_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i1496_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_shr271_i1613_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2__26_i1496_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp296_i1627_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_182to183_bb2_cmp299_i1628_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_or295_i1626_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_lor_ext_i1632_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i1636_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_or295_i1626_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1632_inputs_ready & (local_bb2_or295_i1626_consumed_0_NO_SHIFT_REG | ~(local_bb2_or295_i1626_stall_in)) & local_bb2_lor_ext_i1632_stall_local);
		local_bb2_lor_ext_i1632_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1632_inputs_ready & (local_bb2_lor_ext_i1632_consumed_0_NO_SHIFT_REG | ~(local_bb2_lor_ext_i1632_stall_in)) & local_bb2_lor_ext_i1632_stall_local);
		local_bb2_reduction_0_i1636_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i1632_inputs_ready & (local_bb2_reduction_0_i1636_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i1636_stall_in)) & local_bb2_lor_ext_i1632_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb2_or295_i1078_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1078_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_or295_i1078_0_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1078_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_or295_i1078_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1078_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1078_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1078_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb2_or295_i1078_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb2_or295_i1078_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb2_or295_i1078_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb2_or295_i1078_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb2_or295_i1078_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb2_or295_i1078),
	.data_out(rnode_183to184_bb2_or295_i1078_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb2_or295_i1078_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb2_or295_i1078_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb2_or295_i1078_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb2_or295_i1078_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb2_or295_i1078_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or295_i1078_stall_in = 1'b0;
assign rnode_183to184_bb2_or295_i1078_0_NO_SHIFT_REG = rnode_183to184_bb2_or295_i1078_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb2_or295_i1078_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_or295_i1078_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb2_var__u151_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u151_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_var__u151_0_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u151_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_var__u151_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u151_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u151_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_var__u151_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb2_var__u151_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb2_var__u151_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb2_var__u151_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb2_var__u151_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb2_var__u151_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb2_var__u151),
	.data_out(rnode_183to184_bb2_var__u151_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb2_var__u151_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb2_var__u151_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb2_var__u151_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb2_var__u151_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb2_var__u151_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u151_stall_in = 1'b0;
assign rnode_183to184_bb2_var__u151_0_NO_SHIFT_REG = rnode_183to184_bb2_var__u151_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb2_var__u151_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_var__u151_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb2_lor_ext_i1084_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1084_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_lor_ext_i1084_0_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1084_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_lor_ext_i1084_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1084_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1084_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1084_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb2_lor_ext_i1084_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb2_lor_ext_i1084_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb2_lor_ext_i1084_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb2_lor_ext_i1084_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb2_lor_ext_i1084_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb2_lor_ext_i1084),
	.data_out(rnode_183to184_bb2_lor_ext_i1084_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb2_lor_ext_i1084_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb2_lor_ext_i1084_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb2_lor_ext_i1084_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb2_lor_ext_i1084_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb2_lor_ext_i1084_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lor_ext_i1084_stall_in = 1'b0;
assign rnode_183to184_bb2_lor_ext_i1084_0_NO_SHIFT_REG = rnode_183to184_bb2_lor_ext_i1084_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb2_lor_ext_i1084_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_lor_ext_i1084_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb2_reduction_0_i1088_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1088_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_reduction_0_i1088_0_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1088_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_reduction_0_i1088_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1088_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1088_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1088_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb2_reduction_0_i1088_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb2_reduction_0_i1088_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb2_reduction_0_i1088_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb2_reduction_0_i1088_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb2_reduction_0_i1088_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i1088),
	.data_out(rnode_183to184_bb2_reduction_0_i1088_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb2_reduction_0_i1088_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb2_reduction_0_i1088_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb2_reduction_0_i1088_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb2_reduction_0_i1088_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb2_reduction_0_i1088_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i1088_stall_in = 1'b0;
assign rnode_183to184_bb2_reduction_0_i1088_0_NO_SHIFT_REG = rnode_183to184_bb2_reduction_0_i1088_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb2_reduction_0_i1088_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_reduction_0_i1088_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb2_or295_i1626_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1626_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_or295_i1626_0_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1626_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_or295_i1626_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1626_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1626_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_or295_i1626_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb2_or295_i1626_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb2_or295_i1626_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb2_or295_i1626_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb2_or295_i1626_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb2_or295_i1626_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb2_or295_i1626),
	.data_out(rnode_183to184_bb2_or295_i1626_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb2_or295_i1626_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb2_or295_i1626_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb2_or295_i1626_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb2_or295_i1626_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb2_or295_i1626_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or295_i1626_stall_in = 1'b0;
assign rnode_183to184_bb2_or295_i1626_0_NO_SHIFT_REG = rnode_183to184_bb2_or295_i1626_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb2_or295_i1626_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_or295_i1626_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb2_lor_ext_i1632_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1632_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_lor_ext_i1632_0_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1632_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_lor_ext_i1632_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1632_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1632_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_lor_ext_i1632_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb2_lor_ext_i1632_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb2_lor_ext_i1632_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb2_lor_ext_i1632_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb2_lor_ext_i1632_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb2_lor_ext_i1632_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb2_lor_ext_i1632),
	.data_out(rnode_183to184_bb2_lor_ext_i1632_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb2_lor_ext_i1632_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb2_lor_ext_i1632_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb2_lor_ext_i1632_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb2_lor_ext_i1632_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb2_lor_ext_i1632_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lor_ext_i1632_stall_in = 1'b0;
assign rnode_183to184_bb2_lor_ext_i1632_0_NO_SHIFT_REG = rnode_183to184_bb2_lor_ext_i1632_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb2_lor_ext_i1632_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_lor_ext_i1632_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_183to184_bb2_reduction_0_i1636_0_valid_out_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1636_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_reduction_0_i1636_0_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1636_0_reg_184_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_183to184_bb2_reduction_0_i1636_0_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1636_0_valid_out_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1636_0_stall_in_reg_184_NO_SHIFT_REG;
 logic rnode_183to184_bb2_reduction_0_i1636_0_stall_out_reg_184_NO_SHIFT_REG;

acl_data_fifo rnode_183to184_bb2_reduction_0_i1636_0_reg_184_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_183to184_bb2_reduction_0_i1636_0_reg_184_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_183to184_bb2_reduction_0_i1636_0_stall_in_reg_184_NO_SHIFT_REG),
	.valid_out(rnode_183to184_bb2_reduction_0_i1636_0_valid_out_reg_184_NO_SHIFT_REG),
	.stall_out(rnode_183to184_bb2_reduction_0_i1636_0_stall_out_reg_184_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i1636),
	.data_out(rnode_183to184_bb2_reduction_0_i1636_0_reg_184_NO_SHIFT_REG)
);

defparam rnode_183to184_bb2_reduction_0_i1636_0_reg_184_fifo.DEPTH = 1;
defparam rnode_183to184_bb2_reduction_0_i1636_0_reg_184_fifo.DATA_WIDTH = 32;
defparam rnode_183to184_bb2_reduction_0_i1636_0_reg_184_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_183to184_bb2_reduction_0_i1636_0_reg_184_fifo.IMPL = "shift_reg";

assign rnode_183to184_bb2_reduction_0_i1636_0_reg_184_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i1636_stall_in = 1'b0;
assign rnode_183to184_bb2_reduction_0_i1636_0_NO_SHIFT_REG = rnode_183to184_bb2_reduction_0_i1636_0_reg_184_NO_SHIFT_REG;
assign rnode_183to184_bb2_reduction_0_i1636_0_stall_in_reg_184_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_reduction_0_i1636_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext314_i1087_stall_local;
wire [31:0] local_bb2_lnot_ext314_i1087;

assign local_bb2_lnot_ext314_i1087 = (rnode_183to184_bb2_var__u151_0_NO_SHIFT_REG ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_1_i1637_stall_local;
wire [31:0] local_bb2_reduction_1_i1637;

assign local_bb2_reduction_1_i1637 = (local_bb2_lnot_ext314_i1635 & rnode_183to184_bb2_lor_ext_i1632_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_1_i1089_stall_local;
wire [31:0] local_bb2_reduction_1_i1089;

assign local_bb2_reduction_1_i1089 = (local_bb2_lnot_ext314_i1087 & rnode_183to184_bb2_lor_ext_i1084_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i1638_stall_local;
wire [31:0] local_bb2_reduction_2_i1638;

assign local_bb2_reduction_2_i1638 = (rnode_183to184_bb2_reduction_0_i1636_0_NO_SHIFT_REG & local_bb2_reduction_1_i1637);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i1090_stall_local;
wire [31:0] local_bb2_reduction_2_i1090;

assign local_bb2_reduction_2_i1090 = (rnode_183to184_bb2_reduction_0_i1088_0_NO_SHIFT_REG & local_bb2_reduction_1_i1089);

// This section implements an unregistered operation.
// 
wire local_bb2_add320_i1639_valid_out;
wire local_bb2_add320_i1639_stall_in;
wire local_bb2_add320_i1639_inputs_ready;
wire local_bb2_add320_i1639_stall_local;
wire [31:0] local_bb2_add320_i1639;

assign local_bb2_add320_i1639_inputs_ready = (rnode_183to184_bb2_or295_i1626_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb2_reduction_0_i1636_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb2_var__u150_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb2_lor_ext_i1632_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add320_i1639 = (local_bb2_reduction_2_i1638 + rnode_183to184_bb2_or295_i1626_0_NO_SHIFT_REG);
assign local_bb2_add320_i1639_valid_out = 1'b1;
assign rnode_183to184_bb2_or295_i1626_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_reduction_0_i1636_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_var__u150_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_lor_ext_i1632_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_add320_i1091_valid_out;
wire local_bb2_add320_i1091_stall_in;
wire local_bb2_add320_i1091_inputs_ready;
wire local_bb2_add320_i1091_stall_local;
wire [31:0] local_bb2_add320_i1091;

assign local_bb2_add320_i1091_inputs_ready = (rnode_183to184_bb2_or295_i1078_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb2_reduction_0_i1088_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb2_var__u151_0_valid_out_NO_SHIFT_REG & rnode_183to184_bb2_lor_ext_i1084_0_valid_out_NO_SHIFT_REG);
assign local_bb2_add320_i1091 = (local_bb2_reduction_2_i1090 + rnode_183to184_bb2_or295_i1078_0_NO_SHIFT_REG);
assign local_bb2_add320_i1091_valid_out = 1'b1;
assign rnode_183to184_bb2_or295_i1078_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_reduction_0_i1088_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_var__u151_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_183to184_bb2_lor_ext_i1084_0_stall_in_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb2_add320_i1639_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i1639_0_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i1639_1_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i1639_2_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i1639_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_valid_out_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_stall_in_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1639_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb2_add320_i1639_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb2_add320_i1639_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb2_add320_i1639_0_stall_in_0_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb2_add320_i1639_0_valid_out_0_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb2_add320_i1639_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(local_bb2_add320_i1639),
	.data_out(rnode_184to185_bb2_add320_i1639_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb2_add320_i1639_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb2_add320_i1639_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb2_add320_i1639_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb2_add320_i1639_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb2_add320_i1639_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add320_i1639_stall_in = 1'b0;
assign rnode_184to185_bb2_add320_i1639_0_stall_in_0_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add320_i1639_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i1639_0_NO_SHIFT_REG = rnode_184to185_bb2_add320_i1639_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb2_add320_i1639_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i1639_1_NO_SHIFT_REG = rnode_184to185_bb2_add320_i1639_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb2_add320_i1639_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i1639_2_NO_SHIFT_REG = rnode_184to185_bb2_add320_i1639_0_reg_185_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_184to185_bb2_add320_i1091_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i1091_0_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i1091_1_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i1091_2_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_reg_185_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_184to185_bb2_add320_i1091_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_valid_out_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_stall_in_0_reg_185_NO_SHIFT_REG;
 logic rnode_184to185_bb2_add320_i1091_0_stall_out_reg_185_NO_SHIFT_REG;

acl_data_fifo rnode_184to185_bb2_add320_i1091_0_reg_185_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_184to185_bb2_add320_i1091_0_reg_185_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_184to185_bb2_add320_i1091_0_stall_in_0_reg_185_NO_SHIFT_REG),
	.valid_out(rnode_184to185_bb2_add320_i1091_0_valid_out_0_reg_185_NO_SHIFT_REG),
	.stall_out(rnode_184to185_bb2_add320_i1091_0_stall_out_reg_185_NO_SHIFT_REG),
	.data_in(local_bb2_add320_i1091),
	.data_out(rnode_184to185_bb2_add320_i1091_0_reg_185_NO_SHIFT_REG)
);

defparam rnode_184to185_bb2_add320_i1091_0_reg_185_fifo.DEPTH = 1;
defparam rnode_184to185_bb2_add320_i1091_0_reg_185_fifo.DATA_WIDTH = 32;
defparam rnode_184to185_bb2_add320_i1091_0_reg_185_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_184to185_bb2_add320_i1091_0_reg_185_fifo.IMPL = "shift_reg";

assign rnode_184to185_bb2_add320_i1091_0_reg_185_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add320_i1091_stall_in = 1'b0;
assign rnode_184to185_bb2_add320_i1091_0_stall_in_0_reg_185_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add320_i1091_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i1091_0_NO_SHIFT_REG = rnode_184to185_bb2_add320_i1091_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb2_add320_i1091_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i1091_1_NO_SHIFT_REG = rnode_184to185_bb2_add320_i1091_0_reg_185_NO_SHIFT_REG;
assign rnode_184to185_bb2_add320_i1091_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i1091_2_NO_SHIFT_REG = rnode_184to185_bb2_add320_i1091_0_reg_185_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and2_i448_stall_local;
wire [31:0] local_bb2_and2_i448;

assign local_bb2_and2_i448 = (rnode_184to185_bb2_add320_i1639_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and12_i453_stall_local;
wire [31:0] local_bb2_and12_i453;

assign local_bb2_and12_i453 = (rnode_184to185_bb2_add320_i1639_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb2_add320_i1639_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i1639_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i1639_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i1639_2_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i1639_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1639_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb2_add320_i1639_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb2_add320_i1639_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb2_add320_i1639_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb2_add320_i1639_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb2_add320_i1639_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_184to185_bb2_add320_i1639_2_NO_SHIFT_REG),
	.data_out(rnode_185to186_bb2_add320_i1639_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb2_add320_i1639_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb2_add320_i1639_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_185to186_bb2_add320_i1639_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb2_add320_i1639_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb2_add320_i1639_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i1639_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i1639_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i1639_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i1639_0_NO_SHIFT_REG = rnode_185to186_bb2_add320_i1639_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb2_add320_i1639_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i1639_1_NO_SHIFT_REG = rnode_185to186_bb2_add320_i1639_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb2_add320_i1639_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i1639_2_NO_SHIFT_REG = rnode_185to186_bb2_add320_i1639_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and2_i52_stall_local;
wire [31:0] local_bb2_and2_i52;

assign local_bb2_and2_i52 = (rnode_184to185_bb2_add320_i1091_0_NO_SHIFT_REG >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and12_i_stall_local;
wire [31:0] local_bb2_and12_i;

assign local_bb2_and12_i = (rnode_184to185_bb2_add320_i1091_1_NO_SHIFT_REG & 32'hFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb2_add320_i1091_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i1091_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i1091_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i1091_2_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_185to186_bb2_add320_i1091_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2_add320_i1091_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb2_add320_i1091_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb2_add320_i1091_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb2_add320_i1091_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb2_add320_i1091_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb2_add320_i1091_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(rnode_184to185_bb2_add320_i1091_2_NO_SHIFT_REG),
	.data_out(rnode_185to186_bb2_add320_i1091_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb2_add320_i1091_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb2_add320_i1091_0_reg_186_fifo.DATA_WIDTH = 32;
defparam rnode_185to186_bb2_add320_i1091_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb2_add320_i1091_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb2_add320_i1091_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_184to185_bb2_add320_i1091_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i1091_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i1091_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i1091_0_NO_SHIFT_REG = rnode_185to186_bb2_add320_i1091_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb2_add320_i1091_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i1091_1_NO_SHIFT_REG = rnode_185to186_bb2_add320_i1091_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb2_add320_i1091_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i1091_2_NO_SHIFT_REG = rnode_185to186_bb2_add320_i1091_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i449_stall_local;
wire [31:0] local_bb2_shr3_i449;

assign local_bb2_shr3_i449 = (local_bb2_and2_i448 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp13_i454_stall_local;
wire local_bb2_cmp13_i454;

assign local_bb2_cmp13_i454 = (local_bb2_and10_i452 > local_bb2_and12_i453);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_add320_i1639_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1639_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_add320_i1639_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1639_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_add320_i1639_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1639_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1639_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1639_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_add320_i1639_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_add320_i1639_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_add320_i1639_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_add320_i1639_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_add320_i1639_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(rnode_185to186_bb2_add320_i1639_2_NO_SHIFT_REG),
	.data_out(rnode_186to187_bb2_add320_i1639_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_add320_i1639_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_add320_i1639_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_add320_i1639_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_add320_i1639_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_add320_i1639_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i1639_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_add320_i1639_0_NO_SHIFT_REG = rnode_186to187_bb2_add320_i1639_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_add320_i1639_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_add320_i1639_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_stall_local;
wire [31:0] local_bb2_shr3_i;

assign local_bb2_shr3_i = (local_bb2_and2_i52 & 32'h7FFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp13_i_stall_local;
wire local_bb2_cmp13_i;

assign local_bb2_cmp13_i = (local_bb2_and10_i > local_bb2_and12_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_add320_i1091_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1091_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_add320_i1091_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1091_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_add320_i1091_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1091_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1091_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_add320_i1091_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_add320_i1091_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_add320_i1091_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_add320_i1091_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_add320_i1091_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_add320_i1091_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(rnode_185to186_bb2_add320_i1091_2_NO_SHIFT_REG),
	.data_out(rnode_186to187_bb2_add320_i1091_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_add320_i1091_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_add320_i1091_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_add320_i1091_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_add320_i1091_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_add320_i1091_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2_add320_i1091_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_add320_i1091_0_NO_SHIFT_REG = rnode_186to187_bb2_add320_i1091_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_add320_i1091_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_add320_i1091_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i450_stall_local;
wire local_bb2_cmp_i450;

assign local_bb2_cmp_i450 = (local_bb2_shr_i447 > local_bb2_shr3_i449);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp8_i451_stall_local;
wire local_bb2_cmp8_i451;

assign local_bb2_cmp8_i451 = (local_bb2_shr_i447 == local_bb2_shr3_i449);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_187to190_bb2_add320_i1639_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1639_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to190_bb2_add320_i1639_0_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1639_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to190_bb2_add320_i1639_0_reg_190_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1639_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1639_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1639_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_187to190_bb2_add320_i1639_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to190_bb2_add320_i1639_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to190_bb2_add320_i1639_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_187to190_bb2_add320_i1639_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_187to190_bb2_add320_i1639_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(rnode_186to187_bb2_add320_i1639_0_NO_SHIFT_REG),
	.data_out(rnode_187to190_bb2_add320_i1639_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_187to190_bb2_add320_i1639_0_reg_190_fifo.DEPTH = 3;
defparam rnode_187to190_bb2_add320_i1639_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_187to190_bb2_add320_i1639_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to190_bb2_add320_i1639_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_187to190_bb2_add320_i1639_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_add320_i1639_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_187to190_bb2_add320_i1639_0_NO_SHIFT_REG = rnode_187to190_bb2_add320_i1639_0_reg_190_NO_SHIFT_REG;
assign rnode_187to190_bb2_add320_i1639_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_187to190_bb2_add320_i1639_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp_i53_stall_local;
wire local_bb2_cmp_i53;

assign local_bb2_cmp_i53 = (local_bb2_shr_i51 > local_bb2_shr3_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp8_i_stall_local;
wire local_bb2_cmp8_i;

assign local_bb2_cmp8_i = (local_bb2_shr_i51 == local_bb2_shr3_i);

// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_187to190_bb2_add320_i1091_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1091_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to190_bb2_add320_i1091_0_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1091_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to190_bb2_add320_i1091_0_reg_190_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1091_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1091_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_187to190_bb2_add320_i1091_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_187to190_bb2_add320_i1091_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to190_bb2_add320_i1091_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to190_bb2_add320_i1091_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_187to190_bb2_add320_i1091_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_187to190_bb2_add320_i1091_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(rnode_186to187_bb2_add320_i1091_0_NO_SHIFT_REG),
	.data_out(rnode_187to190_bb2_add320_i1091_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_187to190_bb2_add320_i1091_0_reg_190_fifo.DEPTH = 3;
defparam rnode_187to190_bb2_add320_i1091_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_187to190_bb2_add320_i1091_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to190_bb2_add320_i1091_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_187to190_bb2_add320_i1091_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_add320_i1091_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_187to190_bb2_add320_i1091_0_NO_SHIFT_REG = rnode_187to190_bb2_add320_i1091_0_reg_190_NO_SHIFT_REG;
assign rnode_187to190_bb2_add320_i1091_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_187to190_bb2_add320_i1091_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2___i455_stall_local;
wire local_bb2___i455;

assign local_bb2___i455 = (local_bb2_cmp8_i451 & local_bb2_cmp13_i454);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_add320_i1639_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1639_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_add320_i1639_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1639_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_add320_i1639_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1639_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1639_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1639_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_add320_i1639_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_add320_i1639_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_add320_i1639_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_add320_i1639_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_add320_i1639_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(rnode_187to190_bb2_add320_i1639_0_NO_SHIFT_REG),
	.data_out(rnode_190to191_bb2_add320_i1639_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_add320_i1639_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_add320_i1639_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_add320_i1639_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_add320_i1639_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_add320_i1639_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_187to190_bb2_add320_i1639_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_add320_i1639_0_NO_SHIFT_REG = rnode_190to191_bb2_add320_i1639_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_add320_i1639_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_add320_i1639_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2___i54_stall_local;
wire local_bb2___i54;

assign local_bb2___i54 = (local_bb2_cmp8_i & local_bb2_cmp13_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_add320_i1091_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1091_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_add320_i1091_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1091_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_add320_i1091_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1091_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1091_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_add320_i1091_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_add320_i1091_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_add320_i1091_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_add320_i1091_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_add320_i1091_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_add320_i1091_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(rnode_187to190_bb2_add320_i1091_0_NO_SHIFT_REG),
	.data_out(rnode_190to191_bb2_add320_i1091_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_add320_i1091_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_add320_i1091_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_add320_i1091_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_add320_i1091_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_add320_i1091_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_187to190_bb2_add320_i1091_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_add320_i1091_0_NO_SHIFT_REG = rnode_190to191_bb2_add320_i1091_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_add320_i1091_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_add320_i1091_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2__21_i456_valid_out;
wire local_bb2__21_i456_stall_in;
wire local_bb2__21_i456_inputs_ready;
wire local_bb2__21_i456_stall_local;
wire local_bb2__21_i456;

assign local_bb2__21_i456_inputs_ready = (rnode_184to185_bb2_add320_i1639_0_valid_out_0_NO_SHIFT_REG & rnode_184to185_bb2_add320_i1639_0_valid_out_1_NO_SHIFT_REG & rnode_184to185_bb2_add321_i_0_valid_out_1_NO_SHIFT_REG & rnode_184to185_bb2_add321_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2__21_i456 = (local_bb2_cmp_i450 | local_bb2___i455);
assign local_bb2__21_i456_valid_out = 1'b1;
assign rnode_184to185_bb2_add320_i1639_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add320_i1639_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add321_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add321_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u154_stall_local;
wire [31:0] local_bb2_var__u154;

assign local_bb2_var__u154 = rnode_190to191_bb2_add320_i1639_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__21_i_valid_out;
wire local_bb2__21_i_stall_in;
wire local_bb2__21_i_inputs_ready;
wire local_bb2__21_i_stall_local;
wire local_bb2__21_i;

assign local_bb2__21_i_inputs_ready = (rnode_184to185_bb2_add320_i1091_0_valid_out_0_NO_SHIFT_REG & rnode_184to185_bb2_add320_i1091_0_valid_out_1_NO_SHIFT_REG & rnode_184to185_bb2_add320_i261_0_valid_out_1_NO_SHIFT_REG & rnode_184to185_bb2_add320_i261_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2__21_i = (local_bb2_cmp_i53 | local_bb2___i54);
assign local_bb2__21_i_valid_out = 1'b1;
assign rnode_184to185_bb2_add320_i1091_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add320_i1091_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add320_i261_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_184to185_bb2_add320_i261_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u155_stall_local;
wire [31:0] local_bb2_var__u155;

assign local_bb2_var__u155 = rnode_190to191_bb2_add320_i1091_0_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb2__21_i456_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i456_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb2__21_i456_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb2__21_i456_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb2__21_i456_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb2__21_i456_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb2__21_i456_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb2__21_i456),
	.data_out(rnode_185to186_bb2__21_i456_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb2__21_i456_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb2__21_i456_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb2__21_i456_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb2__21_i456_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb2__21_i456_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__21_i456_stall_in = 1'b0;
assign rnode_185to186_bb2__21_i456_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2__21_i456_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2__21_i456_0_NO_SHIFT_REG = rnode_185to186_bb2__21_i456_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb2__21_i456_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2__21_i456_1_NO_SHIFT_REG = rnode_185to186_bb2__21_i456_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_c0_exi1_stall_local;
wire [159:0] local_bb2_c0_exi1;

assign local_bb2_c0_exi1[31:0] = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
assign local_bb2_c0_exi1[63:32] = local_bb2_var__u154;
assign local_bb2_c0_exi1[159:64] = 96'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_185to186_bb2__21_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_1_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_reg_186_inputs_ready_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_valid_out_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_stall_in_0_reg_186_NO_SHIFT_REG;
 logic rnode_185to186_bb2__21_i_0_stall_out_reg_186_NO_SHIFT_REG;

acl_data_fifo rnode_185to186_bb2__21_i_0_reg_186_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_185to186_bb2__21_i_0_reg_186_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_185to186_bb2__21_i_0_stall_in_0_reg_186_NO_SHIFT_REG),
	.valid_out(rnode_185to186_bb2__21_i_0_valid_out_0_reg_186_NO_SHIFT_REG),
	.stall_out(rnode_185to186_bb2__21_i_0_stall_out_reg_186_NO_SHIFT_REG),
	.data_in(local_bb2__21_i),
	.data_out(rnode_185to186_bb2__21_i_0_reg_186_NO_SHIFT_REG)
);

defparam rnode_185to186_bb2__21_i_0_reg_186_fifo.DEPTH = 1;
defparam rnode_185to186_bb2__21_i_0_reg_186_fifo.DATA_WIDTH = 1;
defparam rnode_185to186_bb2__21_i_0_reg_186_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_185to186_bb2__21_i_0_reg_186_fifo.IMPL = "shift_reg";

assign rnode_185to186_bb2__21_i_0_reg_186_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__21_i_stall_in = 1'b0;
assign rnode_185to186_bb2__21_i_0_stall_in_0_reg_186_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2__21_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2__21_i_0_NO_SHIFT_REG = rnode_185to186_bb2__21_i_0_reg_186_NO_SHIFT_REG;
assign rnode_185to186_bb2__21_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_185to186_bb2__21_i_1_NO_SHIFT_REG = rnode_185to186_bb2__21_i_0_reg_186_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2__22_i457_stall_local;
wire [31:0] local_bb2__22_i457;

assign local_bb2__22_i457 = (rnode_185to186_bb2__21_i456_0_NO_SHIFT_REG ? rnode_185to186_bb2_add320_i1639_0_NO_SHIFT_REG : rnode_185to186_bb2_add321_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2__23_i458_stall_local;
wire [31:0] local_bb2__23_i458;

assign local_bb2__23_i458 = (rnode_185to186_bb2__21_i456_1_NO_SHIFT_REG ? rnode_185to186_bb2_add321_i_1_NO_SHIFT_REG : rnode_185to186_bb2_add320_i1639_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_c0_exi2_stall_local;
wire [159:0] local_bb2_c0_exi2;

assign local_bb2_c0_exi2[63:0] = local_bb2_c0_exi1[63:0];
assign local_bb2_c0_exi2[95:64] = local_bb2_var__u155;
assign local_bb2_c0_exi2[159:96] = local_bb2_c0_exi1[159:96];

// This section implements an unregistered operation.
// 
wire local_bb2__22_i_stall_local;
wire [31:0] local_bb2__22_i;

assign local_bb2__22_i = (rnode_185to186_bb2__21_i_0_NO_SHIFT_REG ? rnode_185to186_bb2_add320_i1091_0_NO_SHIFT_REG : rnode_185to186_bb2_add320_i261_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2__23_i_stall_local;
wire [31:0] local_bb2__23_i;

assign local_bb2__23_i = (rnode_185to186_bb2__21_i_1_NO_SHIFT_REG ? rnode_185to186_bb2_add320_i261_1_NO_SHIFT_REG : rnode_185to186_bb2_add320_i1091_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shr18_i461_stall_local;
wire [31:0] local_bb2_shr18_i461;

assign local_bb2_shr18_i461 = (local_bb2__22_i457 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i459_stall_local;
wire [31:0] local_bb2_shr16_i459;

assign local_bb2_shr16_i459 = (local_bb2__23_i458 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shr18_i_stall_local;
wire [31:0] local_bb2_shr18_i;

assign local_bb2_shr18_i = (local_bb2__22_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_shr16_i_stall_local;
wire [31:0] local_bb2_shr16_i;

assign local_bb2_shr16_i = (local_bb2__23_i >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and19_i462_stall_local;
wire [31:0] local_bb2_and19_i462;

assign local_bb2_and19_i462 = (local_bb2_shr18_i461 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i491_stall_local;
wire [31:0] local_bb2_sub_i491;

assign local_bb2_sub_i491 = (local_bb2_shr16_i459 - local_bb2_shr18_i461);

// This section implements an unregistered operation.
// 
wire local_bb2_and19_i_stall_local;
wire [31:0] local_bb2_and19_i;

assign local_bb2_and19_i = (local_bb2_shr18_i & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_sub_i63_stall_local;
wire [31:0] local_bb2_sub_i63;

assign local_bb2_sub_i63 = (local_bb2_shr16_i - local_bb2_shr18_i);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot23_i466_stall_local;
wire local_bb2_lnot23_i466;

assign local_bb2_lnot23_i466 = (local_bb2_and19_i462 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp27_i468_stall_local;
wire local_bb2_cmp27_i468;

assign local_bb2_cmp27_i468 = (local_bb2_and19_i462 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and68_i492_stall_local;
wire [31:0] local_bb2_and68_i492;

assign local_bb2_and68_i492 = (local_bb2_sub_i491 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot23_i_stall_local;
wire local_bb2_lnot23_i;

assign local_bb2_lnot23_i = (local_bb2_and19_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp27_i_stall_local;
wire local_bb2_cmp27_i;

assign local_bb2_cmp27_i = (local_bb2_and19_i == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and68_i_stall_local;
wire [31:0] local_bb2_and68_i;

assign local_bb2_and68_i = (local_bb2_sub_i63 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp69_i493_stall_local;
wire local_bb2_cmp69_i493;

assign local_bb2_cmp69_i493 = (local_bb2_and68_i492 > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp69_i_stall_local;
wire local_bb2_cmp69_i;

assign local_bb2_cmp69_i = (local_bb2_and68_i > 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_align_0_i494_stall_local;
wire [31:0] local_bb2_align_0_i494;

assign local_bb2_align_0_i494 = (local_bb2_cmp69_i493 ? 32'h1F : local_bb2_and68_i492);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i_valid_out_1;
wire local_bb2__22_i_stall_in_1;
 reg local_bb2__22_i_consumed_1_NO_SHIFT_REG;
wire local_bb2__23_i_valid_out_1;
wire local_bb2__23_i_stall_in_1;
 reg local_bb2__23_i_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr16_i_valid_out_1;
wire local_bb2_shr16_i_stall_in_1;
 reg local_bb2_shr16_i_consumed_1_NO_SHIFT_REG;
wire local_bb2_lnot23_i_valid_out;
wire local_bb2_lnot23_i_stall_in;
 reg local_bb2_lnot23_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp27_i_valid_out;
wire local_bb2_cmp27_i_stall_in;
 reg local_bb2_cmp27_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i_valid_out;
wire local_bb2_align_0_i_stall_in;
 reg local_bb2_align_0_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_align_0_i_inputs_ready;
wire local_bb2_align_0_i_stall_local;
wire [31:0] local_bb2_align_0_i;

assign local_bb2_align_0_i_inputs_ready = (rnode_185to186_bb2__21_i_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb2_add320_i1091_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb2_add320_i261_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb2__21_i_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb2_add320_i1091_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb2_add320_i261_0_valid_out_1_NO_SHIFT_REG);
assign local_bb2_align_0_i = (local_bb2_cmp69_i ? 32'h1F : local_bb2_and68_i);
assign local_bb2__22_i_valid_out_1 = 1'b1;
assign local_bb2__23_i_valid_out_1 = 1'b1;
assign local_bb2_shr16_i_valid_out_1 = 1'b1;
assign local_bb2_lnot23_i_valid_out = 1'b1;
assign local_bb2_cmp27_i_valid_out = 1'b1;
assign local_bb2_align_0_i_valid_out = 1'b1;
assign rnode_185to186_bb2__21_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i1091_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i261_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2__21_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i1091_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i261_0_stall_in_1_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__22_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__23_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr16_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lnot23_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp27_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_align_0_i_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__22_i_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i_inputs_ready & (local_bb2__22_i_consumed_1_NO_SHIFT_REG | ~(local_bb2__22_i_stall_in_1)) & local_bb2_align_0_i_stall_local);
		local_bb2__23_i_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i_inputs_ready & (local_bb2__23_i_consumed_1_NO_SHIFT_REG | ~(local_bb2__23_i_stall_in_1)) & local_bb2_align_0_i_stall_local);
		local_bb2_shr16_i_consumed_1_NO_SHIFT_REG <= (local_bb2_align_0_i_inputs_ready & (local_bb2_shr16_i_consumed_1_NO_SHIFT_REG | ~(local_bb2_shr16_i_stall_in_1)) & local_bb2_align_0_i_stall_local);
		local_bb2_lnot23_i_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i_inputs_ready & (local_bb2_lnot23_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_lnot23_i_stall_in)) & local_bb2_align_0_i_stall_local);
		local_bb2_cmp27_i_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i_inputs_ready & (local_bb2_cmp27_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp27_i_stall_in)) & local_bb2_align_0_i_stall_local);
		local_bb2_align_0_i_consumed_0_NO_SHIFT_REG <= (local_bb2_align_0_i_inputs_ready & (local_bb2_align_0_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_align_0_i_stall_in)) & local_bb2_align_0_i_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_and93_i502_stall_local;
wire [31:0] local_bb2_and93_i502;

assign local_bb2_and93_i502 = (local_bb2_align_0_i494 & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb2_and95_i504_stall_local;
wire [31:0] local_bb2_and95_i504;

assign local_bb2_and95_i504 = (local_bb2_align_0_i494 & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and115_i520_stall_local;
wire [31:0] local_bb2_and115_i520;

assign local_bb2_and115_i520 = (local_bb2_align_0_i494 & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_and130_i526_stall_local;
wire [31:0] local_bb2_and130_i526;

assign local_bb2_and130_i526 = (local_bb2_align_0_i494 & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2__22_i457_valid_out_1;
wire local_bb2__22_i457_stall_in_1;
 reg local_bb2__22_i457_consumed_1_NO_SHIFT_REG;
wire local_bb2__23_i458_valid_out_1;
wire local_bb2__23_i458_stall_in_1;
 reg local_bb2__23_i458_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr16_i459_valid_out_1;
wire local_bb2_shr16_i459_stall_in_1;
 reg local_bb2_shr16_i459_consumed_1_NO_SHIFT_REG;
wire local_bb2_lnot23_i466_valid_out;
wire local_bb2_lnot23_i466_stall_in;
 reg local_bb2_lnot23_i466_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp27_i468_valid_out;
wire local_bb2_cmp27_i468_stall_in;
 reg local_bb2_cmp27_i468_consumed_0_NO_SHIFT_REG;
wire local_bb2_and93_i502_valid_out;
wire local_bb2_and93_i502_stall_in;
 reg local_bb2_and93_i502_consumed_0_NO_SHIFT_REG;
wire local_bb2_and95_i504_valid_out;
wire local_bb2_and95_i504_stall_in;
 reg local_bb2_and95_i504_consumed_0_NO_SHIFT_REG;
wire local_bb2_and115_i520_valid_out;
wire local_bb2_and115_i520_stall_in;
 reg local_bb2_and115_i520_consumed_0_NO_SHIFT_REG;
wire local_bb2_and130_i526_valid_out;
wire local_bb2_and130_i526_stall_in;
 reg local_bb2_and130_i526_consumed_0_NO_SHIFT_REG;
wire local_bb2_and149_i531_valid_out;
wire local_bb2_and149_i531_stall_in;
 reg local_bb2_and149_i531_consumed_0_NO_SHIFT_REG;
wire local_bb2_and149_i531_inputs_ready;
wire local_bb2_and149_i531_stall_local;
wire [31:0] local_bb2_and149_i531;

assign local_bb2_and149_i531_inputs_ready = (rnode_185to186_bb2__21_i456_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb2_add320_i1639_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb2_add321_i_0_valid_out_0_NO_SHIFT_REG & rnode_185to186_bb2__21_i456_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb2_add320_i1639_0_valid_out_1_NO_SHIFT_REG & rnode_185to186_bb2_add321_i_0_valid_out_1_NO_SHIFT_REG);
assign local_bb2_and149_i531 = (local_bb2_align_0_i494 & 32'h3);
assign local_bb2__22_i457_valid_out_1 = 1'b1;
assign local_bb2__23_i458_valid_out_1 = 1'b1;
assign local_bb2_shr16_i459_valid_out_1 = 1'b1;
assign local_bb2_lnot23_i466_valid_out = 1'b1;
assign local_bb2_cmp27_i468_valid_out = 1'b1;
assign local_bb2_and93_i502_valid_out = 1'b1;
assign local_bb2_and95_i504_valid_out = 1'b1;
assign local_bb2_and115_i520_valid_out = 1'b1;
assign local_bb2_and130_i526_valid_out = 1'b1;
assign local_bb2_and149_i531_valid_out = 1'b1;
assign rnode_185to186_bb2__21_i456_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i1639_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add321_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2__21_i456_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add320_i1639_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_185to186_bb2_add321_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2__22_i457_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__23_i458_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr16_i459_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lnot23_i466_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp27_i468_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and93_i502_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and95_i504_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and115_i520_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and130_i526_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and149_i531_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2__22_i457_consumed_1_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2__22_i457_consumed_1_NO_SHIFT_REG | ~(local_bb2__22_i457_stall_in_1)) & local_bb2_and149_i531_stall_local);
		local_bb2__23_i458_consumed_1_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2__23_i458_consumed_1_NO_SHIFT_REG | ~(local_bb2__23_i458_stall_in_1)) & local_bb2_and149_i531_stall_local);
		local_bb2_shr16_i459_consumed_1_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2_shr16_i459_consumed_1_NO_SHIFT_REG | ~(local_bb2_shr16_i459_stall_in_1)) & local_bb2_and149_i531_stall_local);
		local_bb2_lnot23_i466_consumed_0_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2_lnot23_i466_consumed_0_NO_SHIFT_REG | ~(local_bb2_lnot23_i466_stall_in)) & local_bb2_and149_i531_stall_local);
		local_bb2_cmp27_i468_consumed_0_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2_cmp27_i468_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp27_i468_stall_in)) & local_bb2_and149_i531_stall_local);
		local_bb2_and93_i502_consumed_0_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2_and93_i502_consumed_0_NO_SHIFT_REG | ~(local_bb2_and93_i502_stall_in)) & local_bb2_and149_i531_stall_local);
		local_bb2_and95_i504_consumed_0_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2_and95_i504_consumed_0_NO_SHIFT_REG | ~(local_bb2_and95_i504_stall_in)) & local_bb2_and149_i531_stall_local);
		local_bb2_and115_i520_consumed_0_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2_and115_i520_consumed_0_NO_SHIFT_REG | ~(local_bb2_and115_i520_stall_in)) & local_bb2_and149_i531_stall_local);
		local_bb2_and130_i526_consumed_0_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2_and130_i526_consumed_0_NO_SHIFT_REG | ~(local_bb2_and130_i526_stall_in)) & local_bb2_and149_i531_stall_local);
		local_bb2_and149_i531_consumed_0_NO_SHIFT_REG <= (local_bb2_and149_i531_inputs_ready & (local_bb2_and149_i531_consumed_0_NO_SHIFT_REG | ~(local_bb2_and149_i531_stall_in)) & local_bb2_and149_i531_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2__22_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__22_i_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__22_i_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__22_i_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2__22_i_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2__22_i_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2__22_i_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2__22_i_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2__22_i_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2__22_i),
	.data_out(rnode_186to187_bb2__22_i_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2__22_i_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2__22_i_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2__22_i_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2__22_i_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2__22_i_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__22_i_stall_in_1 = 1'b0;
assign rnode_186to187_bb2__22_i_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__22_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__22_i_0_NO_SHIFT_REG = rnode_186to187_bb2__22_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2__22_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__22_i_1_NO_SHIFT_REG = rnode_186to187_bb2__22_i_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2__23_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__23_i_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__23_i_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__23_i_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__23_i_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2__23_i_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2__23_i_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2__23_i_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2__23_i_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2__23_i_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2__23_i),
	.data_out(rnode_186to187_bb2__23_i_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2__23_i_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2__23_i_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2__23_i_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2__23_i_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2__23_i_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__23_i_stall_in_1 = 1'b0;
assign rnode_186to187_bb2__23_i_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__23_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__23_i_0_NO_SHIFT_REG = rnode_186to187_bb2__23_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2__23_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__23_i_1_NO_SHIFT_REG = rnode_186to187_bb2__23_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2__23_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__23_i_2_NO_SHIFT_REG = rnode_186to187_bb2__23_i_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_shr16_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_shr16_i_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_shr16_i_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_shr16_i_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_shr16_i_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_shr16_i_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_shr16_i_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_shr16_i_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_shr16_i_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_shr16_i),
	.data_out(rnode_186to187_bb2_shr16_i_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_shr16_i_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_shr16_i_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_shr16_i_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_shr16_i_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_shr16_i_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr16_i_stall_in_1 = 1'b0;
assign rnode_186to187_bb2_shr16_i_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_shr16_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_shr16_i_0_NO_SHIFT_REG = rnode_186to187_bb2_shr16_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_shr16_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_shr16_i_1_NO_SHIFT_REG = rnode_186to187_bb2_shr16_i_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_lnot23_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_lnot23_i_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_lnot23_i_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_lnot23_i_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_lnot23_i_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_lnot23_i_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_lnot23_i),
	.data_out(rnode_186to187_bb2_lnot23_i_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_lnot23_i_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_lnot23_i_0_reg_187_fifo.DATA_WIDTH = 1;
defparam rnode_186to187_bb2_lnot23_i_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_lnot23_i_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_lnot23_i_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lnot23_i_stall_in = 1'b0;
assign rnode_186to187_bb2_lnot23_i_0_NO_SHIFT_REG = rnode_186to187_bb2_lnot23_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_lnot23_i_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_lnot23_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_cmp27_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_cmp27_i_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_cmp27_i_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_cmp27_i_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_cmp27_i_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_cmp27_i_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_cmp27_i),
	.data_out(rnode_186to187_bb2_cmp27_i_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_cmp27_i_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_cmp27_i_0_reg_187_fifo.DATA_WIDTH = 1;
defparam rnode_186to187_bb2_cmp27_i_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_cmp27_i_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_cmp27_i_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp27_i_stall_in = 1'b0;
assign rnode_186to187_bb2_cmp27_i_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_cmp27_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_cmp27_i_0_NO_SHIFT_REG = rnode_186to187_bb2_cmp27_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_cmp27_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_cmp27_i_1_NO_SHIFT_REG = rnode_186to187_bb2_cmp27_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_cmp27_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_cmp27_i_2_NO_SHIFT_REG = rnode_186to187_bb2_cmp27_i_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_align_0_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_align_0_i_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_align_0_i_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_align_0_i_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_align_0_i_3_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_valid_out_4_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_stall_in_4_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_align_0_i_4_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_align_0_i_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_align_0_i_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_align_0_i_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_align_0_i_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_align_0_i_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_align_0_i_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_align_0_i_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_align_0_i),
	.data_out(rnode_186to187_bb2_align_0_i_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_align_0_i_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_align_0_i_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_align_0_i_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_align_0_i_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_align_0_i_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_align_0_i_stall_in = 1'b0;
assign rnode_186to187_bb2_align_0_i_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_align_0_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_align_0_i_0_NO_SHIFT_REG = rnode_186to187_bb2_align_0_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_align_0_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_align_0_i_1_NO_SHIFT_REG = rnode_186to187_bb2_align_0_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_align_0_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_align_0_i_2_NO_SHIFT_REG = rnode_186to187_bb2_align_0_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_align_0_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_align_0_i_3_NO_SHIFT_REG = rnode_186to187_bb2_align_0_i_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_align_0_i_0_valid_out_4_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_align_0_i_4_NO_SHIFT_REG = rnode_186to187_bb2_align_0_i_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2__22_i457_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i457_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__22_i457_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i457_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i457_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__22_i457_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i457_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__22_i457_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i457_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i457_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__22_i457_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2__22_i457_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2__22_i457_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2__22_i457_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2__22_i457_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2__22_i457_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2__22_i457),
	.data_out(rnode_186to187_bb2__22_i457_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2__22_i457_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2__22_i457_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2__22_i457_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2__22_i457_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2__22_i457_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__22_i457_stall_in_1 = 1'b0;
assign rnode_186to187_bb2__22_i457_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__22_i457_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__22_i457_0_NO_SHIFT_REG = rnode_186to187_bb2__22_i457_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2__22_i457_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__22_i457_1_NO_SHIFT_REG = rnode_186to187_bb2__22_i457_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2__23_i458_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__23_i458_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__23_i458_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__23_i458_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2__23_i458_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2__23_i458_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2__23_i458_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2__23_i458_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2__23_i458_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2__23_i458_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2__23_i458_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2__23_i458),
	.data_out(rnode_186to187_bb2__23_i458_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2__23_i458_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2__23_i458_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2__23_i458_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2__23_i458_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2__23_i458_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__23_i458_stall_in_1 = 1'b0;
assign rnode_186to187_bb2__23_i458_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__23_i458_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__23_i458_0_NO_SHIFT_REG = rnode_186to187_bb2__23_i458_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2__23_i458_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__23_i458_1_NO_SHIFT_REG = rnode_186to187_bb2__23_i458_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2__23_i458_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2__23_i458_2_NO_SHIFT_REG = rnode_186to187_bb2__23_i458_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_shr16_i459_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i459_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_shr16_i459_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i459_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i459_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_shr16_i459_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i459_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_shr16_i459_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i459_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i459_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_shr16_i459_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_shr16_i459_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_shr16_i459_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_shr16_i459_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_shr16_i459_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_shr16_i459_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_shr16_i459),
	.data_out(rnode_186to187_bb2_shr16_i459_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_shr16_i459_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_shr16_i459_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_shr16_i459_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_shr16_i459_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_shr16_i459_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr16_i459_stall_in_1 = 1'b0;
assign rnode_186to187_bb2_shr16_i459_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_shr16_i459_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_shr16_i459_0_NO_SHIFT_REG = rnode_186to187_bb2_shr16_i459_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_shr16_i459_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_shr16_i459_1_NO_SHIFT_REG = rnode_186to187_bb2_shr16_i459_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_lnot23_i466_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i466_0_stall_in_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i466_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i466_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i466_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i466_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i466_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_lnot23_i466_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_lnot23_i466_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_lnot23_i466_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_lnot23_i466_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_lnot23_i466_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_lnot23_i466_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_lnot23_i466),
	.data_out(rnode_186to187_bb2_lnot23_i466_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_lnot23_i466_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_lnot23_i466_0_reg_187_fifo.DATA_WIDTH = 1;
defparam rnode_186to187_bb2_lnot23_i466_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_lnot23_i466_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_lnot23_i466_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lnot23_i466_stall_in = 1'b0;
assign rnode_186to187_bb2_lnot23_i466_0_NO_SHIFT_REG = rnode_186to187_bb2_lnot23_i466_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_lnot23_i466_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_lnot23_i466_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_cmp27_i468_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_cmp27_i468_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_cmp27_i468_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_cmp27_i468_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_cmp27_i468_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_cmp27_i468_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_cmp27_i468_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_cmp27_i468),
	.data_out(rnode_186to187_bb2_cmp27_i468_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_cmp27_i468_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_cmp27_i468_0_reg_187_fifo.DATA_WIDTH = 1;
defparam rnode_186to187_bb2_cmp27_i468_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_cmp27_i468_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_cmp27_i468_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp27_i468_stall_in = 1'b0;
assign rnode_186to187_bb2_cmp27_i468_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_cmp27_i468_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_cmp27_i468_0_NO_SHIFT_REG = rnode_186to187_bb2_cmp27_i468_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_cmp27_i468_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_cmp27_i468_1_NO_SHIFT_REG = rnode_186to187_bb2_cmp27_i468_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_cmp27_i468_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_cmp27_i468_2_NO_SHIFT_REG = rnode_186to187_bb2_cmp27_i468_0_reg_187_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_and93_i502_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and93_i502_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and93_i502_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and93_i502_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and93_i502_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and93_i502_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and93_i502_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and93_i502_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_and93_i502_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_and93_i502_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_and93_i502_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_and93_i502_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_and93_i502_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_and93_i502),
	.data_out(rnode_186to187_bb2_and93_i502_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_and93_i502_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_and93_i502_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_and93_i502_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_and93_i502_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_and93_i502_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and93_i502_stall_in = 1'b0;
assign rnode_186to187_bb2_and93_i502_0_NO_SHIFT_REG = rnode_186to187_bb2_and93_i502_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_and93_i502_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and93_i502_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_and95_i504_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and95_i504_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and95_i504_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and95_i504_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and95_i504_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and95_i504_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and95_i504_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and95_i504_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_and95_i504_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_and95_i504_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_and95_i504_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_and95_i504_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_and95_i504_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_and95_i504),
	.data_out(rnode_186to187_bb2_and95_i504_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_and95_i504_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_and95_i504_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_and95_i504_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_and95_i504_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_and95_i504_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and95_i504_stall_in = 1'b0;
assign rnode_186to187_bb2_and95_i504_0_NO_SHIFT_REG = rnode_186to187_bb2_and95_i504_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_and95_i504_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and95_i504_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_and115_i520_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and115_i520_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and115_i520_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and115_i520_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and115_i520_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and115_i520_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and115_i520_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and115_i520_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_and115_i520_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_and115_i520_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_and115_i520_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_and115_i520_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_and115_i520_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_and115_i520),
	.data_out(rnode_186to187_bb2_and115_i520_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_and115_i520_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_and115_i520_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_and115_i520_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_and115_i520_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_and115_i520_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and115_i520_stall_in = 1'b0;
assign rnode_186to187_bb2_and115_i520_0_NO_SHIFT_REG = rnode_186to187_bb2_and115_i520_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_and115_i520_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and115_i520_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_and130_i526_0_valid_out_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and130_i526_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and130_i526_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and130_i526_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and130_i526_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and130_i526_0_valid_out_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and130_i526_0_stall_in_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and130_i526_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_and130_i526_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_and130_i526_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_and130_i526_0_stall_in_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_and130_i526_0_valid_out_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_and130_i526_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_and130_i526),
	.data_out(rnode_186to187_bb2_and130_i526_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_and130_i526_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_and130_i526_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_and130_i526_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_and130_i526_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_and130_i526_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and130_i526_stall_in = 1'b0;
assign rnode_186to187_bb2_and130_i526_0_NO_SHIFT_REG = rnode_186to187_bb2_and130_i526_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_and130_i526_0_stall_in_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and130_i526_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_186to187_bb2_and149_i531_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and149_i531_0_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and149_i531_1_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and149_i531_2_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_reg_187_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_186to187_bb2_and149_i531_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_valid_out_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_stall_in_0_reg_187_NO_SHIFT_REG;
 logic rnode_186to187_bb2_and149_i531_0_stall_out_reg_187_NO_SHIFT_REG;

acl_data_fifo rnode_186to187_bb2_and149_i531_0_reg_187_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_186to187_bb2_and149_i531_0_reg_187_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_186to187_bb2_and149_i531_0_stall_in_0_reg_187_NO_SHIFT_REG),
	.valid_out(rnode_186to187_bb2_and149_i531_0_valid_out_0_reg_187_NO_SHIFT_REG),
	.stall_out(rnode_186to187_bb2_and149_i531_0_stall_out_reg_187_NO_SHIFT_REG),
	.data_in(local_bb2_and149_i531),
	.data_out(rnode_186to187_bb2_and149_i531_0_reg_187_NO_SHIFT_REG)
);

defparam rnode_186to187_bb2_and149_i531_0_reg_187_fifo.DEPTH = 1;
defparam rnode_186to187_bb2_and149_i531_0_reg_187_fifo.DATA_WIDTH = 32;
defparam rnode_186to187_bb2_and149_i531_0_reg_187_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_186to187_bb2_and149_i531_0_reg_187_fifo.IMPL = "shift_reg";

assign rnode_186to187_bb2_and149_i531_0_reg_187_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and149_i531_stall_in = 1'b0;
assign rnode_186to187_bb2_and149_i531_0_stall_in_0_reg_187_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and149_i531_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_and149_i531_0_NO_SHIFT_REG = rnode_186to187_bb2_and149_i531_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_and149_i531_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_and149_i531_1_NO_SHIFT_REG = rnode_186to187_bb2_and149_i531_0_reg_187_NO_SHIFT_REG;
assign rnode_186to187_bb2_and149_i531_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_and149_i531_2_NO_SHIFT_REG = rnode_186to187_bb2_and149_i531_0_reg_187_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and21_i_stall_local;
wire [31:0] local_bb2_and21_i;

assign local_bb2_and21_i = (rnode_186to187_bb2__22_i_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and20_i_stall_local;
wire [31:0] local_bb2_and20_i;

assign local_bb2_and20_i = (rnode_186to187_bb2__23_i_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and35_i_valid_out;
wire local_bb2_and35_i_stall_in;
wire local_bb2_and35_i_inputs_ready;
wire local_bb2_and35_i_stall_local;
wire [31:0] local_bb2_and35_i;

assign local_bb2_and35_i_inputs_ready = rnode_186to187_bb2__23_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and35_i = (rnode_186to187_bb2__23_i_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb2_and35_i_valid_out = 1'b1;
assign rnode_186to187_bb2__23_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i57_stall_local;
wire [31:0] local_bb2_xor_i57;

assign local_bb2_xor_i57 = (rnode_186to187_bb2__23_i_2_NO_SHIFT_REG ^ rnode_186to187_bb2__22_i_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and17_i_stall_local;
wire [31:0] local_bb2_and17_i;

assign local_bb2_and17_i = (rnode_186to187_bb2_shr16_i_0_NO_SHIFT_REG & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_187to189_bb2_shr16_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to189_bb2_shr16_i_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to189_bb2_shr16_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_187to189_bb2_shr16_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to189_bb2_shr16_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to189_bb2_shr16_i_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_187to189_bb2_shr16_i_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_187to189_bb2_shr16_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(rnode_186to187_bb2_shr16_i_1_NO_SHIFT_REG),
	.data_out(rnode_187to189_bb2_shr16_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_187to189_bb2_shr16_i_0_reg_189_fifo.DEPTH = 2;
defparam rnode_187to189_bb2_shr16_i_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_187to189_bb2_shr16_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to189_bb2_shr16_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_187to189_bb2_shr16_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_shr16_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_shr16_i_0_NO_SHIFT_REG = rnode_187to189_bb2_shr16_i_0_reg_189_NO_SHIFT_REG;
assign rnode_187to189_bb2_shr16_i_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_shr16_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and93_i_stall_local;
wire [31:0] local_bb2_and93_i;

assign local_bb2_and93_i = (rnode_186to187_bb2_align_0_i_0_NO_SHIFT_REG & 32'h1C);

// This section implements an unregistered operation.
// 
wire local_bb2_and95_i_stall_local;
wire [31:0] local_bb2_and95_i;

assign local_bb2_and95_i = (rnode_186to187_bb2_align_0_i_1_NO_SHIFT_REG & 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_and115_i_stall_local;
wire [31:0] local_bb2_and115_i;

assign local_bb2_and115_i = (rnode_186to187_bb2_align_0_i_2_NO_SHIFT_REG & 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_and130_i_stall_local;
wire [31:0] local_bb2_and130_i;

assign local_bb2_and130_i = (rnode_186to187_bb2_align_0_i_3_NO_SHIFT_REG & 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and149_i_stall_local;
wire [31:0] local_bb2_and149_i;

assign local_bb2_and149_i = (rnode_186to187_bb2_align_0_i_4_NO_SHIFT_REG & 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and21_i464_stall_local;
wire [31:0] local_bb2_and21_i464;

assign local_bb2_and21_i464 = (rnode_186to187_bb2__22_i457_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and20_i463_stall_local;
wire [31:0] local_bb2_and20_i463;

assign local_bb2_and20_i463 = (rnode_186to187_bb2__23_i458_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and35_i469_valid_out;
wire local_bb2_and35_i469_stall_in;
wire local_bb2_and35_i469_inputs_ready;
wire local_bb2_and35_i469_stall_local;
wire [31:0] local_bb2_and35_i469;

assign local_bb2_and35_i469_inputs_ready = rnode_186to187_bb2__23_i458_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and35_i469 = (rnode_186to187_bb2__23_i458_1_NO_SHIFT_REG & 32'h80000000);
assign local_bb2_and35_i469_valid_out = 1'b1;
assign rnode_186to187_bb2__23_i458_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_xor_i470_stall_local;
wire [31:0] local_bb2_xor_i470;

assign local_bb2_xor_i470 = (rnode_186to187_bb2__23_i458_2_NO_SHIFT_REG ^ rnode_186to187_bb2__22_i457_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and17_i460_stall_local;
wire [31:0] local_bb2_and17_i460;

assign local_bb2_and17_i460 = (rnode_186to187_bb2_shr16_i459_0_NO_SHIFT_REG & 32'hFF);

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_187to189_bb2_shr16_i459_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i459_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to189_bb2_shr16_i459_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i459_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to189_bb2_shr16_i459_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i459_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i459_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_shr16_i459_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_187to189_bb2_shr16_i459_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to189_bb2_shr16_i459_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to189_bb2_shr16_i459_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_187to189_bb2_shr16_i459_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_187to189_bb2_shr16_i459_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(rnode_186to187_bb2_shr16_i459_1_NO_SHIFT_REG),
	.data_out(rnode_187to189_bb2_shr16_i459_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_187to189_bb2_shr16_i459_0_reg_189_fifo.DEPTH = 2;
defparam rnode_187to189_bb2_shr16_i459_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_187to189_bb2_shr16_i459_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to189_bb2_shr16_i459_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_187to189_bb2_shr16_i459_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_186to187_bb2_shr16_i459_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_shr16_i459_0_NO_SHIFT_REG = rnode_187to189_bb2_shr16_i459_0_reg_189_NO_SHIFT_REG;
assign rnode_187to189_bb2_shr16_i459_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_shr16_i459_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp96_i505_stall_local;
wire local_bb2_cmp96_i505;

assign local_bb2_cmp96_i505 = (rnode_186to187_bb2_and95_i504_0_NO_SHIFT_REG == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp116_i521_stall_local;
wire local_bb2_cmp116_i521;

assign local_bb2_cmp116_i521 = (rnode_186to187_bb2_and115_i520_0_NO_SHIFT_REG == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp131_not_i528_stall_local;
wire local_bb2_cmp131_not_i528;

assign local_bb2_cmp131_not_i528 = (rnode_186to187_bb2_and130_i526_0_NO_SHIFT_REG != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_Pivot20_i533_stall_local;
wire local_bb2_Pivot20_i533;

assign local_bb2_Pivot20_i533 = (rnode_186to187_bb2_and149_i531_1_NO_SHIFT_REG < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_SwitchLeaf_i534_stall_local;
wire local_bb2_SwitchLeaf_i534;

assign local_bb2_SwitchLeaf_i534 = (rnode_186to187_bb2_and149_i531_2_NO_SHIFT_REG == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot33_not_i_stall_local;
wire local_bb2_lnot33_not_i;

assign local_bb2_lnot33_not_i = (local_bb2_and21_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or64_i_stall_local;
wire [31:0] local_bb2_or64_i;

assign local_bb2_or64_i = (local_bb2_and21_i << 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_i_stall_local;
wire local_bb2_lnot30_i;

assign local_bb2_lnot30_i = (local_bb2_and20_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i59_stall_local;
wire [31:0] local_bb2_or_i59;

assign local_bb2_or_i59 = (local_bb2_and20_i << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb2_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_and35_i_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_and35_i_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb2_and35_i_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb2_and35_i_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb2_and35_i_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb2_and35_i_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb2_and35_i_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb2_and35_i),
	.data_out(rnode_187to188_bb2_and35_i_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb2_and35_i_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb2_and35_i_0_reg_188_fifo.DATA_WIDTH = 32;
defparam rnode_187to188_bb2_and35_i_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb2_and35_i_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb2_and35_i_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and35_i_stall_in = 1'b0;
assign rnode_187to188_bb2_and35_i_0_NO_SHIFT_REG = rnode_187to188_bb2_and35_i_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_and35_i_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb2_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i_stall_local;
wire local_bb2_cmp37_i;

assign local_bb2_cmp37_i = ($signed(local_bb2_xor_i57) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_xor_lobit_i_stall_local;
wire [31:0] local_bb2_xor_lobit_i;

assign local_bb2_xor_lobit_i = ($signed(local_bb2_xor_i57) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and36_lobit_i_stall_local;
wire [31:0] local_bb2_and36_lobit_i;

assign local_bb2_and36_lobit_i = (local_bb2_xor_i57 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i55_stall_local;
wire local_bb2_lnot_i55;

assign local_bb2_lnot_i55 = (local_bb2_and17_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_i56_stall_local;
wire local_bb2_cmp25_i56;

assign local_bb2_cmp25_i56 = (local_bb2_and17_i == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp96_i_stall_local;
wire local_bb2_cmp96_i;

assign local_bb2_cmp96_i = (local_bb2_and95_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp116_i_stall_local;
wire local_bb2_cmp116_i;

assign local_bb2_cmp116_i = (local_bb2_and115_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp131_not_i_stall_local;
wire local_bb2_cmp131_not_i;

assign local_bb2_cmp131_not_i = (local_bb2_and130_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_Pivot20_i_stall_local;
wire local_bb2_Pivot20_i;

assign local_bb2_Pivot20_i = (local_bb2_and149_i < 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_SwitchLeaf_i_stall_local;
wire local_bb2_SwitchLeaf_i;

assign local_bb2_SwitchLeaf_i = (local_bb2_and149_i == 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot33_not_i475_stall_local;
wire local_bb2_lnot33_not_i475;

assign local_bb2_lnot33_not_i475 = (local_bb2_and21_i464 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or64_i488_stall_local;
wire [31:0] local_bb2_or64_i488;

assign local_bb2_or64_i488 = (local_bb2_and21_i464 << 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_i473_stall_local;
wire local_bb2_lnot30_i473;

assign local_bb2_lnot30_i473 = (local_bb2_and20_i463 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i485_stall_local;
wire [31:0] local_bb2_or_i485;

assign local_bb2_or_i485 = (local_bb2_and20_i463 << 32'h3);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb2_and35_i469_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i469_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_and35_i469_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i469_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_and35_i469_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i469_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i469_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_and35_i469_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb2_and35_i469_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb2_and35_i469_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb2_and35_i469_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb2_and35_i469_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb2_and35_i469_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb2_and35_i469),
	.data_out(rnode_187to188_bb2_and35_i469_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb2_and35_i469_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb2_and35_i469_0_reg_188_fifo.DATA_WIDTH = 32;
defparam rnode_187to188_bb2_and35_i469_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb2_and35_i469_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb2_and35_i469_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and35_i469_stall_in = 1'b0;
assign rnode_187to188_bb2_and35_i469_0_NO_SHIFT_REG = rnode_187to188_bb2_and35_i469_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_and35_i469_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb2_and35_i469_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i471_stall_local;
wire local_bb2_cmp37_i471;

assign local_bb2_cmp37_i471 = ($signed(local_bb2_xor_i470) < $signed(32'h0));

// This section implements an unregistered operation.
// 
wire local_bb2_xor_lobit_i544_stall_local;
wire [31:0] local_bb2_xor_lobit_i544;

assign local_bb2_xor_lobit_i544 = ($signed(local_bb2_xor_i470) >>> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and36_lobit_i546_stall_local;
wire [31:0] local_bb2_and36_lobit_i546;

assign local_bb2_and36_lobit_i546 = (local_bb2_xor_i470 >> 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_i465_stall_local;
wire local_bb2_lnot_i465;

assign local_bb2_lnot_i465 = (local_bb2_and17_i460 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_i467_stall_local;
wire local_bb2_cmp25_i467;

assign local_bb2_cmp25_i467 = (local_bb2_and17_i460 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_i_stall_local;
wire local_bb2_brmerge_not_i;

assign local_bb2_brmerge_not_i = (rnode_186to187_bb2_cmp27_i_0_NO_SHIFT_REG & local_bb2_lnot33_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_shl65_i_stall_local;
wire [31:0] local_bb2_shl65_i;

assign local_bb2_shl65_i = (local_bb2_or64_i | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_not_i_stall_local;
wire local_bb2_lnot30_not_i;

assign local_bb2_lnot30_not_i = (local_bb2_lnot30_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i60_stall_local;
wire [31:0] local_bb2_shl_i60;

assign local_bb2_shl_i60 = (local_bb2_or_i59 | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and35_i_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and35_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_and35_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_and35_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_and35_i_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_and35_i_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_and35_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(rnode_187to188_bb2_and35_i_0_NO_SHIFT_REG),
	.data_out(rnode_188to189_bb2_and35_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_and35_i_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_and35_i_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2_and35_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_and35_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_and35_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and35_i_0_NO_SHIFT_REG = rnode_188to189_bb2_and35_i_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and35_i_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_not_i_stall_local;
wire local_bb2_cmp25_not_i;

assign local_bb2_cmp25_not_i = (local_bb2_cmp25_i56 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u156_stall_local;
wire local_bb2_var__u156;

assign local_bb2_var__u156 = (local_bb2_cmp25_i56 | rnode_186to187_bb2_cmp27_i_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_i476_stall_local;
wire local_bb2_brmerge_not_i476;

assign local_bb2_brmerge_not_i476 = (rnode_186to187_bb2_cmp27_i468_0_NO_SHIFT_REG & local_bb2_lnot33_not_i475);

// This section implements an unregistered operation.
// 
wire local_bb2_shl65_i489_stall_local;
wire [31:0] local_bb2_shl65_i489;

assign local_bb2_shl65_i489 = (local_bb2_or64_i488 | 32'h4000000);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot30_not_i477_stall_local;
wire local_bb2_lnot30_not_i477;

assign local_bb2_lnot30_not_i477 = (local_bb2_lnot30_i473 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_shl_i486_stall_local;
wire [31:0] local_bb2_shl_i486;

assign local_bb2_shl_i486 = (local_bb2_or_i485 | 32'h4000000);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_and35_i469_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i469_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and35_i469_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i469_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and35_i469_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i469_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i469_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and35_i469_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_and35_i469_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_and35_i469_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_and35_i469_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_and35_i469_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_and35_i469_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(rnode_187to188_bb2_and35_i469_0_NO_SHIFT_REG),
	.data_out(rnode_188to189_bb2_and35_i469_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_and35_i469_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_and35_i469_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2_and35_i469_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_and35_i469_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_and35_i469_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_and35_i469_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and35_i469_0_NO_SHIFT_REG = rnode_188to189_bb2_and35_i469_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and35_i469_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and35_i469_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp25_not_i472_stall_local;
wire local_bb2_cmp25_not_i472;

assign local_bb2_cmp25_not_i472 = (local_bb2_cmp25_i467 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u157_stall_local;
wire local_bb2_var__u157;

assign local_bb2_var__u157 = (local_bb2_cmp25_i467 | rnode_186to187_bb2_cmp27_i468_2_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_not_i_stall_local;
wire local_bb2_brmerge_not_not_i;

assign local_bb2_brmerge_not_not_i = (local_bb2_brmerge_not_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i62_stall_local;
wire [31:0] local_bb2__28_i62;

assign local_bb2__28_i62 = (rnode_186to187_bb2_lnot23_i_0_NO_SHIFT_REG ? 32'h0 : local_bb2_shl65_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_not_i_stall_local;
wire local_bb2_or_cond_not_i;

assign local_bb2_or_cond_not_i = (local_bb2_cmp25_i56 & local_bb2_lnot30_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i61_stall_local;
wire [31:0] local_bb2__27_i61;

assign local_bb2__27_i61 = (local_bb2_lnot_i55 ? 32'h0 : local_bb2_shl_i60);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_and35_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_and35_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_and35_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_and35_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_and35_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_and35_i_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_and35_i_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_and35_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(rnode_188to189_bb2_and35_i_0_NO_SHIFT_REG),
	.data_out(rnode_189to190_bb2_and35_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_and35_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_and35_i_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_189to190_bb2_and35_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_and35_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_and35_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_and35_i_0_NO_SHIFT_REG = rnode_189to190_bb2_and35_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_and35_i_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_and35_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_i_stall_local;
wire local_bb2_or_cond_i;

assign local_bb2_or_cond_i = (local_bb2_lnot30_i | local_bb2_cmp25_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge_not_not_i480_stall_local;
wire local_bb2_brmerge_not_not_i480;

assign local_bb2_brmerge_not_not_i480 = (local_bb2_brmerge_not_i476 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__28_i490_stall_local;
wire [31:0] local_bb2__28_i490;

assign local_bb2__28_i490 = (rnode_186to187_bb2_lnot23_i466_0_NO_SHIFT_REG ? 32'h0 : local_bb2_shl65_i489);

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_not_i478_stall_local;
wire local_bb2_or_cond_not_i478;

assign local_bb2_or_cond_not_i478 = (local_bb2_cmp25_i467 & local_bb2_lnot30_not_i477);

// This section implements an unregistered operation.
// 
wire local_bb2__27_i487_stall_local;
wire [31:0] local_bb2__27_i487;

assign local_bb2__27_i487 = (local_bb2_lnot_i465 ? 32'h0 : local_bb2_shl_i486);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_and35_i469_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i469_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_and35_i469_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i469_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_and35_i469_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i469_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i469_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and35_i469_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_and35_i469_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_and35_i469_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_and35_i469_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_and35_i469_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_and35_i469_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(rnode_188to189_bb2_and35_i469_0_NO_SHIFT_REG),
	.data_out(rnode_189to190_bb2_and35_i469_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_and35_i469_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_and35_i469_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_189to190_bb2_and35_i469_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_and35_i469_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_and35_i469_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_and35_i469_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_and35_i469_0_NO_SHIFT_REG = rnode_189to190_bb2_and35_i469_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_and35_i469_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_and35_i469_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_or_cond_i474_stall_local;
wire local_bb2_or_cond_i474;

assign local_bb2_or_cond_i474 = (local_bb2_lnot30_i473 | local_bb2_cmp25_not_i472);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_7_i_stall_local;
wire local_bb2_reduction_7_i;

assign local_bb2_reduction_7_i = (local_bb2_cmp25_i56 & local_bb2_brmerge_not_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_i_stall_local;
wire [31:0] local_bb2_and72_i;

assign local_bb2_and72_i = (local_bb2__28_i62 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i64_stall_local;
wire [31:0] local_bb2_and75_i64;

assign local_bb2_and75_i64 = (local_bb2__28_i62 & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb2_and78_i_stall_local;
wire [31:0] local_bb2_and78_i;

assign local_bb2_and78_i = (local_bb2__28_i62 & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb2_shr94_i_stall_local;
wire [31:0] local_bb2_shr94_i;

assign local_bb2_shr94_i = (local_bb2__28_i62 >> local_bb2_and93_i);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i65_stall_local;
wire [31:0] local_bb2_and90_i65;

assign local_bb2_and90_i65 = (local_bb2__28_i62 & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and87_i_stall_local;
wire [31:0] local_bb2_and87_i;

assign local_bb2_and87_i = (local_bb2__28_i62 & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb2_and84_i_stall_local;
wire [31:0] local_bb2_and84_i;

assign local_bb2_and84_i = (local_bb2__28_i62 & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u158_stall_local;
wire [31:0] local_bb2_var__u158;

assign local_bb2_var__u158 = (local_bb2__28_i62 & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i58_stall_local;
wire local_bb2__24_i58;

assign local_bb2__24_i58 = (local_bb2_or_cond_not_i | local_bb2_brmerge_not_i);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i74_stall_local;
wire [31:0] local_bb2_add_i74;

assign local_bb2_add_i74 = (local_bb2__27_i61 | local_bb2_and36_lobit_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_8_i_stall_local;
wire local_bb2_reduction_8_i;

assign local_bb2_reduction_8_i = (rnode_186to187_bb2_cmp27_i_1_NO_SHIFT_REG & local_bb2_or_cond_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_7_i481_stall_local;
wire local_bb2_reduction_7_i481;

assign local_bb2_reduction_7_i481 = (local_bb2_cmp25_i467 & local_bb2_brmerge_not_not_i480);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_i495_stall_local;
wire [31:0] local_bb2_and72_i495;

assign local_bb2_and72_i495 = (local_bb2__28_i490 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and75_i498_stall_local;
wire [31:0] local_bb2_and75_i498;

assign local_bb2_and75_i498 = (local_bb2__28_i490 & 32'hF0);

// This section implements an unregistered operation.
// 
wire local_bb2_and78_i500_stall_local;
wire [31:0] local_bb2_and78_i500;

assign local_bb2_and78_i500 = (local_bb2__28_i490 & 32'hF00);

// This section implements an unregistered operation.
// 
wire local_bb2_shr94_i503_stall_local;
wire [31:0] local_bb2_shr94_i503;

assign local_bb2_shr94_i503 = (local_bb2__28_i490 >> rnode_186to187_bb2_and93_i502_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_and90_i506_stall_local;
wire [31:0] local_bb2_and90_i506;

assign local_bb2_and90_i506 = (local_bb2__28_i490 & 32'h7000000);

// This section implements an unregistered operation.
// 
wire local_bb2_and87_i507_stall_local;
wire [31:0] local_bb2_and87_i507;

assign local_bb2_and87_i507 = (local_bb2__28_i490 & 32'hF00000);

// This section implements an unregistered operation.
// 
wire local_bb2_and84_i508_stall_local;
wire [31:0] local_bb2_and84_i508;

assign local_bb2_and84_i508 = (local_bb2__28_i490 & 32'hF0000);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u159_stall_local;
wire [31:0] local_bb2_var__u159;

assign local_bb2_var__u159 = (local_bb2__28_i490 & 32'hFFF8);

// This section implements an unregistered operation.
// 
wire local_bb2__24_i479_stall_local;
wire local_bb2__24_i479;

assign local_bb2__24_i479 = (local_bb2_or_cond_not_i478 | local_bb2_brmerge_not_i476);

// This section implements an unregistered operation.
// 
wire local_bb2_add_i547_stall_local;
wire [31:0] local_bb2_add_i547;

assign local_bb2_add_i547 = (local_bb2__27_i487 | local_bb2_and36_lobit_i546);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_8_i482_stall_local;
wire local_bb2_reduction_8_i482;

assign local_bb2_reduction_8_i482 = (rnode_186to187_bb2_cmp27_i468_1_NO_SHIFT_REG & local_bb2_or_cond_i474);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_tr_i_stall_local;
wire [7:0] local_bb2_and72_tr_i;

assign local_bb2_and72_tr_i = local_bb2_and72_i[7:0];

// This section implements an unregistered operation.
// 
wire local_bb2_cmp76_i_stall_local;
wire local_bb2_cmp76_i;

assign local_bb2_cmp76_i = (local_bb2_and75_i64 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp79_i_stall_local;
wire local_bb2_cmp79_i;

assign local_bb2_cmp79_i = (local_bb2_and78_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_and142_i_stall_local;
wire [31:0] local_bb2_and142_i;

assign local_bb2_and142_i = (local_bb2_shr94_i >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr150_i_stall_local;
wire [31:0] local_bb2_shr150_i;

assign local_bb2_shr150_i = (local_bb2_shr94_i >> local_bb2_and149_i);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u160_stall_local;
wire [31:0] local_bb2_var__u160;

assign local_bb2_var__u160 = (local_bb2_shr94_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and146_i_stall_local;
wire [31:0] local_bb2_and146_i;

assign local_bb2_and146_i = (local_bb2_shr94_i >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i66_stall_local;
wire local_bb2_cmp91_i66;

assign local_bb2_cmp91_i66 = (local_bb2_and90_i65 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp88_i_stall_local;
wire local_bb2_cmp88_i;

assign local_bb2_cmp88_i = (local_bb2_and87_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp85_i_stall_local;
wire local_bb2_cmp85_i;

assign local_bb2_cmp85_i = (local_bb2_and84_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u161_stall_local;
wire local_bb2_var__u161;

assign local_bb2_var__u161 = (local_bb2_var__u158 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_9_i_stall_local;
wire local_bb2_reduction_9_i;

assign local_bb2_reduction_9_i = (local_bb2_reduction_7_i & local_bb2_reduction_8_i);

// This section implements an unregistered operation.
// 
wire local_bb2_and72_tr_i496_stall_local;
wire [7:0] local_bb2_and72_tr_i496;

assign local_bb2_and72_tr_i496 = local_bb2_and72_i495[7:0];

// This section implements an unregistered operation.
// 
wire local_bb2_cmp76_i499_stall_local;
wire local_bb2_cmp76_i499;

assign local_bb2_cmp76_i499 = (local_bb2_and75_i498 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp79_i501_stall_local;
wire local_bb2_cmp79_i501;

assign local_bb2_cmp79_i501 = (local_bb2_and78_i500 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_and142_i530_stall_local;
wire [31:0] local_bb2_and142_i530;

assign local_bb2_and142_i530 = (local_bb2_shr94_i503 >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_shr150_i532_stall_local;
wire [31:0] local_bb2_shr150_i532;

assign local_bb2_shr150_i532 = (local_bb2_shr94_i503 >> rnode_186to187_bb2_and149_i531_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u162_stall_local;
wire [31:0] local_bb2_var__u162;

assign local_bb2_var__u162 = (local_bb2_shr94_i503 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and146_i535_stall_local;
wire [31:0] local_bb2_and146_i535;

assign local_bb2_and146_i535 = (local_bb2_shr94_i503 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp91_i509_stall_local;
wire local_bb2_cmp91_i509;

assign local_bb2_cmp91_i509 = (local_bb2_and90_i506 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp88_i510_stall_local;
wire local_bb2_cmp88_i510;

assign local_bb2_cmp88_i510 = (local_bb2_and87_i507 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp85_i511_stall_local;
wire local_bb2_cmp85_i511;

assign local_bb2_cmp85_i511 = (local_bb2_and84_i508 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u163_stall_local;
wire local_bb2_var__u163;

assign local_bb2_var__u163 = (local_bb2_var__u159 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_9_i483_stall_local;
wire local_bb2_reduction_9_i483;

assign local_bb2_reduction_9_i483 = (local_bb2_reduction_7_i481 & local_bb2_reduction_8_i482);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool74_i_stall_local;
wire [7:0] local_bb2_frombool74_i;

assign local_bb2_frombool74_i = (local_bb2_and72_tr_i & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u164_stall_local;
wire [31:0] local_bb2_var__u164;

assign local_bb2_var__u164 = (local_bb2_and146_i | local_bb2_shr94_i);

// This section implements an unregistered operation.
// 
wire local_bb2__31_v_i_stall_local;
wire local_bb2__31_v_i;

assign local_bb2__31_v_i = (local_bb2_cmp96_i ? local_bb2_cmp79_i : local_bb2_cmp91_i66);

// This section implements an unregistered operation.
// 
wire local_bb2__30_v_i_stall_local;
wire local_bb2__30_v_i;

assign local_bb2__30_v_i = (local_bb2_cmp96_i ? local_bb2_cmp76_i : local_bb2_cmp88_i);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool109_i_stall_local;
wire [7:0] local_bb2_frombool109_i;

assign local_bb2_frombool109_i[7:1] = 7'h0;
assign local_bb2_frombool109_i[0] = local_bb2_cmp85_i;

// This section implements an unregistered operation.
// 
wire local_bb2_or107_i_stall_local;
wire [31:0] local_bb2_or107_i;

assign local_bb2_or107_i[31:1] = 31'h0;
assign local_bb2_or107_i[0] = local_bb2_var__u161;

// This section implements an unregistered operation.
// 
wire local_bb2__26_i_stall_local;
wire local_bb2__26_i;

assign local_bb2__26_i = (local_bb2_reduction_9_i ? local_bb2_cmp37_i : local_bb2__24_i58);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool74_i497_stall_local;
wire [7:0] local_bb2_frombool74_i497;

assign local_bb2_frombool74_i497 = (local_bb2_and72_tr_i496 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u165_stall_local;
wire [31:0] local_bb2_var__u165;

assign local_bb2_var__u165 = (local_bb2_and146_i535 | local_bb2_shr94_i503);

// This section implements an unregistered operation.
// 
wire local_bb2__31_v_i517_stall_local;
wire local_bb2__31_v_i517;

assign local_bb2__31_v_i517 = (local_bb2_cmp96_i505 ? local_bb2_cmp79_i501 : local_bb2_cmp91_i509);

// This section implements an unregistered operation.
// 
wire local_bb2__30_v_i515_stall_local;
wire local_bb2__30_v_i515;

assign local_bb2__30_v_i515 = (local_bb2_cmp96_i505 ? local_bb2_cmp76_i499 : local_bb2_cmp88_i510);

// This section implements an unregistered operation.
// 
wire local_bb2_frombool109_i513_stall_local;
wire [7:0] local_bb2_frombool109_i513;

assign local_bb2_frombool109_i513[7:1] = 7'h0;
assign local_bb2_frombool109_i513[0] = local_bb2_cmp85_i511;

// This section implements an unregistered operation.
// 
wire local_bb2_or107_i512_stall_local;
wire [31:0] local_bb2_or107_i512;

assign local_bb2_or107_i512[31:1] = 31'h0;
assign local_bb2_or107_i512[0] = local_bb2_var__u163;

// This section implements an unregistered operation.
// 
wire local_bb2__26_i484_stall_local;
wire local_bb2__26_i484;

assign local_bb2__26_i484 = (local_bb2_reduction_9_i483 ? local_bb2_cmp37_i471 : local_bb2__24_i479);

// This section implements an unregistered operation.
// 
wire local_bb2_or1596_i_stall_local;
wire [31:0] local_bb2_or1596_i;

assign local_bb2_or1596_i = (local_bb2_var__u164 | local_bb2_and142_i);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i68_stall_local;
wire [7:0] local_bb2__31_i68;

assign local_bb2__31_i68[7:1] = 7'h0;
assign local_bb2__31_i68[0] = local_bb2__31_v_i;

// This section implements an unregistered operation.
// 
wire local_bb2__30_i_stall_local;
wire [7:0] local_bb2__30_i;

assign local_bb2__30_i[7:1] = 7'h0;
assign local_bb2__30_i[0] = local_bb2__30_v_i;

// This section implements an unregistered operation.
// 
wire local_bb2__29_i67_stall_local;
wire [7:0] local_bb2__29_i67;

assign local_bb2__29_i67 = (local_bb2_cmp96_i ? local_bb2_frombool74_i : local_bb2_frombool109_i);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i69_stall_local;
wire [31:0] local_bb2__32_i69;

assign local_bb2__32_i69 = (local_bb2_cmp96_i ? 32'h0 : local_bb2_or107_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or1596_i536_stall_local;
wire [31:0] local_bb2_or1596_i536;

assign local_bb2_or1596_i536 = (local_bb2_var__u165 | local_bb2_and142_i530);

// This section implements an unregistered operation.
// 
wire local_bb2__31_i518_stall_local;
wire [7:0] local_bb2__31_i518;

assign local_bb2__31_i518[7:1] = 7'h0;
assign local_bb2__31_i518[0] = local_bb2__31_v_i517;

// This section implements an unregistered operation.
// 
wire local_bb2__30_i516_stall_local;
wire [7:0] local_bb2__30_i516;

assign local_bb2__30_i516[7:1] = 7'h0;
assign local_bb2__30_i516[0] = local_bb2__30_v_i515;

// This section implements an unregistered operation.
// 
wire local_bb2__29_i514_stall_local;
wire [7:0] local_bb2__29_i514;

assign local_bb2__29_i514 = (local_bb2_cmp96_i505 ? local_bb2_frombool74_i497 : local_bb2_frombool109_i513);

// This section implements an unregistered operation.
// 
wire local_bb2__32_i519_stall_local;
wire [31:0] local_bb2__32_i519;

assign local_bb2__32_i519 = (local_bb2_cmp96_i505 ? 32'h0 : local_bb2_or107_i512);

// This section implements an unregistered operation.
// 
wire local_bb2_or162_i_stall_local;
wire [31:0] local_bb2_or162_i;

assign local_bb2_or162_i = (local_bb2_or1596_i & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or1237_i_stall_local;
wire [7:0] local_bb2_or1237_i;

assign local_bb2_or1237_i = (local_bb2__30_i | local_bb2__29_i67);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i70_stall_local;
wire [7:0] local_bb2__33_i70;

assign local_bb2__33_i70 = (local_bb2_cmp116_i ? local_bb2__29_i67 : local_bb2__31_i68);

// This section implements an unregistered operation.
// 
wire local_bb2_or162_i537_stall_local;
wire [31:0] local_bb2_or162_i537;

assign local_bb2_or162_i537 = (local_bb2_or1596_i536 & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or1237_i522_stall_local;
wire [7:0] local_bb2_or1237_i522;

assign local_bb2_or1237_i522 = (local_bb2__30_i516 | local_bb2__29_i514);

// This section implements an unregistered operation.
// 
wire local_bb2__33_i524_stall_local;
wire [7:0] local_bb2__33_i524;

assign local_bb2__33_i524 = (local_bb2_cmp116_i521 ? local_bb2__29_i514 : local_bb2__31_i518);

// This section implements an unregistered operation.
// 
wire local_bb2__37_v_i_stall_local;
wire [31:0] local_bb2__37_v_i;

assign local_bb2__37_v_i = (local_bb2_Pivot20_i ? 32'h0 : local_bb2_or162_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or123_i_stall_local;
wire [31:0] local_bb2_or123_i;

assign local_bb2_or123_i[31:8] = 24'h0;
assign local_bb2_or123_i[7:0] = local_bb2_or1237_i;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u166_stall_local;
wire [7:0] local_bb2_var__u166;

assign local_bb2_var__u166 = (local_bb2__33_i70 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__37_v_i538_stall_local;
wire [31:0] local_bb2__37_v_i538;

assign local_bb2__37_v_i538 = (local_bb2_Pivot20_i533 ? 32'h0 : local_bb2_or162_i537);

// This section implements an unregistered operation.
// 
wire local_bb2_or123_i523_stall_local;
wire [31:0] local_bb2_or123_i523;

assign local_bb2_or123_i523[31:8] = 24'h0;
assign local_bb2_or123_i523[7:0] = local_bb2_or1237_i522;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u167_stall_local;
wire [7:0] local_bb2_var__u167;

assign local_bb2_var__u167 = (local_bb2__33_i524 & 8'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__39_v_i_stall_local;
wire [31:0] local_bb2__39_v_i;

assign local_bb2__39_v_i = (local_bb2_SwitchLeaf_i ? local_bb2_var__u160 : local_bb2__37_v_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or124_i_stall_local;
wire [31:0] local_bb2_or124_i;

assign local_bb2_or124_i = (local_bb2_cmp116_i ? 32'h0 : local_bb2_or123_i);

// This section implements an unregistered operation.
// 
wire local_bb2_conv135_i_stall_local;
wire [31:0] local_bb2_conv135_i;

assign local_bb2_conv135_i[31:8] = 24'h0;
assign local_bb2_conv135_i[7:0] = local_bb2_var__u166;

// This section implements an unregistered operation.
// 
wire local_bb2__39_v_i539_stall_local;
wire [31:0] local_bb2__39_v_i539;

assign local_bb2__39_v_i539 = (local_bb2_SwitchLeaf_i534 ? local_bb2_var__u162 : local_bb2__37_v_i538);

// This section implements an unregistered operation.
// 
wire local_bb2_or124_i525_stall_local;
wire [31:0] local_bb2_or124_i525;

assign local_bb2_or124_i525 = (local_bb2_cmp116_i521 ? 32'h0 : local_bb2_or123_i523);

// This section implements an unregistered operation.
// 
wire local_bb2_conv135_i527_stall_local;
wire [31:0] local_bb2_conv135_i527;

assign local_bb2_conv135_i527[31:8] = 24'h0;
assign local_bb2_conv135_i527[7:0] = local_bb2_var__u167;

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i71_stall_local;
wire [31:0] local_bb2_reduction_3_i71;

assign local_bb2_reduction_3_i71 = (local_bb2__32_i69 | local_bb2_or124_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or136_i_stall_local;
wire [31:0] local_bb2_or136_i;

assign local_bb2_or136_i = (local_bb2_cmp131_not_i ? local_bb2_conv135_i : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_3_i540_stall_local;
wire [31:0] local_bb2_reduction_3_i540;

assign local_bb2_reduction_3_i540 = (local_bb2__32_i519 | local_bb2_or124_i525);

// This section implements an unregistered operation.
// 
wire local_bb2_or136_i529_stall_local;
wire [31:0] local_bb2_or136_i529;

assign local_bb2_or136_i529 = (local_bb2_cmp131_not_i528 ? local_bb2_conv135_i527 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i72_stall_local;
wire [31:0] local_bb2_reduction_5_i72;

assign local_bb2_reduction_5_i72 = (local_bb2_shr150_i | local_bb2_reduction_3_i71);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_4_i_stall_local;
wire [31:0] local_bb2_reduction_4_i;

assign local_bb2_reduction_4_i = (local_bb2_or136_i | local_bb2__39_v_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_5_i542_stall_local;
wire [31:0] local_bb2_reduction_5_i542;

assign local_bb2_reduction_5_i542 = (local_bb2_shr150_i532 | local_bb2_reduction_3_i540);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_4_i541_stall_local;
wire [31:0] local_bb2_reduction_4_i541;

assign local_bb2_reduction_4_i541 = (local_bb2_or136_i529 | local_bb2__39_v_i539);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i73_stall_local;
wire [31:0] local_bb2_reduction_6_i73;

assign local_bb2_reduction_6_i73 = (local_bb2_reduction_4_i | local_bb2_reduction_5_i72);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_6_i543_stall_local;
wire [31:0] local_bb2_reduction_6_i543;

assign local_bb2_reduction_6_i543 = (local_bb2_reduction_4_i541 | local_bb2_reduction_5_i542);

// This section implements an unregistered operation.
// 
wire local_bb2_xor188_i_stall_local;
wire [31:0] local_bb2_xor188_i;

assign local_bb2_xor188_i = (local_bb2_reduction_6_i73 ^ local_bb2_xor_lobit_i);

// This section implements an unregistered operation.
// 
wire local_bb2_xor188_i545_stall_local;
wire [31:0] local_bb2_xor188_i545;

assign local_bb2_xor188_i545 = (local_bb2_reduction_6_i543 ^ local_bb2_xor_lobit_i544);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i_valid_out_1;
wire local_bb2_cmp37_i_stall_in_1;
 reg local_bb2_cmp37_i_consumed_1_NO_SHIFT_REG;
wire local_bb2__26_i_valid_out;
wire local_bb2__26_i_stall_in;
 reg local_bb2__26_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i_valid_out;
wire local_bb2_add192_i_stall_in;
 reg local_bb2_add192_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_and17_i_valid_out_2;
wire local_bb2_and17_i_stall_in_2;
 reg local_bb2_and17_i_consumed_2_NO_SHIFT_REG;
wire local_bb2_var__u156_valid_out;
wire local_bb2_var__u156_stall_in;
 reg local_bb2_var__u156_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i_inputs_ready;
wire local_bb2_add192_i_stall_local;
wire [31:0] local_bb2_add192_i;

assign local_bb2_add192_i_inputs_ready = (rnode_186to187_bb2__22_i_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_cmp27_i_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_lnot23_i_0_valid_out_NO_SHIFT_REG & rnode_186to187_bb2__23_i_0_valid_out_2_NO_SHIFT_REG & rnode_186to187_bb2__22_i_0_valid_out_1_NO_SHIFT_REG & rnode_186to187_bb2__23_i_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_cmp27_i_0_valid_out_1_NO_SHIFT_REG & rnode_186to187_bb2_shr16_i_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_cmp27_i_0_valid_out_2_NO_SHIFT_REG & rnode_186to187_bb2_align_0_i_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_align_0_i_0_valid_out_4_NO_SHIFT_REG & rnode_186to187_bb2_align_0_i_0_valid_out_1_NO_SHIFT_REG & rnode_186to187_bb2_align_0_i_0_valid_out_2_NO_SHIFT_REG & rnode_186to187_bb2_align_0_i_0_valid_out_3_NO_SHIFT_REG);
assign local_bb2_add192_i = (local_bb2_add_i74 + local_bb2_xor188_i);
assign local_bb2_cmp37_i_valid_out_1 = 1'b1;
assign local_bb2__26_i_valid_out = 1'b1;
assign local_bb2_add192_i_valid_out = 1'b1;
assign local_bb2_and17_i_valid_out_2 = 1'b1;
assign local_bb2_var__u156_valid_out = 1'b1;
assign rnode_186to187_bb2__22_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_cmp27_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_lnot23_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__23_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__22_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__23_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_cmp27_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_shr16_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_cmp27_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_align_0_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_align_0_i_0_stall_in_4_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_align_0_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_align_0_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_align_0_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp37_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__26_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add192_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and17_i_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u156_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp37_i_consumed_1_NO_SHIFT_REG <= (local_bb2_add192_i_inputs_ready & (local_bb2_cmp37_i_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp37_i_stall_in_1)) & local_bb2_add192_i_stall_local);
		local_bb2__26_i_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i_inputs_ready & (local_bb2__26_i_consumed_0_NO_SHIFT_REG | ~(local_bb2__26_i_stall_in)) & local_bb2_add192_i_stall_local);
		local_bb2_add192_i_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i_inputs_ready & (local_bb2_add192_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_add192_i_stall_in)) & local_bb2_add192_i_stall_local);
		local_bb2_and17_i_consumed_2_NO_SHIFT_REG <= (local_bb2_add192_i_inputs_ready & (local_bb2_and17_i_consumed_2_NO_SHIFT_REG | ~(local_bb2_and17_i_stall_in_2)) & local_bb2_add192_i_stall_local);
		local_bb2_var__u156_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i_inputs_ready & (local_bb2_var__u156_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u156_stall_in)) & local_bb2_add192_i_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp37_i471_valid_out_1;
wire local_bb2_cmp37_i471_stall_in_1;
 reg local_bb2_cmp37_i471_consumed_1_NO_SHIFT_REG;
wire local_bb2__26_i484_valid_out;
wire local_bb2__26_i484_stall_in;
 reg local_bb2__26_i484_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i548_valid_out;
wire local_bb2_add192_i548_stall_in;
 reg local_bb2_add192_i548_consumed_0_NO_SHIFT_REG;
wire local_bb2_and17_i460_valid_out_2;
wire local_bb2_and17_i460_stall_in_2;
 reg local_bb2_and17_i460_consumed_2_NO_SHIFT_REG;
wire local_bb2_var__u157_valid_out;
wire local_bb2_var__u157_stall_in;
 reg local_bb2_var__u157_consumed_0_NO_SHIFT_REG;
wire local_bb2_add192_i548_inputs_ready;
wire local_bb2_add192_i548_stall_local;
wire [31:0] local_bb2_add192_i548;

assign local_bb2_add192_i548_inputs_ready = (rnode_186to187_bb2__22_i457_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_cmp27_i468_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_lnot23_i466_0_valid_out_NO_SHIFT_REG & rnode_186to187_bb2_and93_i502_0_valid_out_NO_SHIFT_REG & rnode_186to187_bb2__23_i458_0_valid_out_2_NO_SHIFT_REG & rnode_186to187_bb2__22_i457_0_valid_out_1_NO_SHIFT_REG & rnode_186to187_bb2__23_i458_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_cmp27_i468_0_valid_out_1_NO_SHIFT_REG & rnode_186to187_bb2_shr16_i459_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_cmp27_i468_0_valid_out_2_NO_SHIFT_REG & rnode_186to187_bb2_and149_i531_0_valid_out_0_NO_SHIFT_REG & rnode_186to187_bb2_and95_i504_0_valid_out_NO_SHIFT_REG & rnode_186to187_bb2_and149_i531_0_valid_out_2_NO_SHIFT_REG & rnode_186to187_bb2_and115_i520_0_valid_out_NO_SHIFT_REG & rnode_186to187_bb2_and130_i526_0_valid_out_NO_SHIFT_REG & rnode_186to187_bb2_and149_i531_0_valid_out_1_NO_SHIFT_REG);
assign local_bb2_add192_i548 = (local_bb2_add_i547 + local_bb2_xor188_i545);
assign local_bb2_cmp37_i471_valid_out_1 = 1'b1;
assign local_bb2__26_i484_valid_out = 1'b1;
assign local_bb2_add192_i548_valid_out = 1'b1;
assign local_bb2_and17_i460_valid_out_2 = 1'b1;
assign local_bb2_var__u157_valid_out = 1'b1;
assign rnode_186to187_bb2__22_i457_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_cmp27_i468_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_lnot23_i466_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and93_i502_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__23_i458_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__22_i457_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2__23_i458_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_cmp27_i468_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_shr16_i459_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_cmp27_i468_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and149_i531_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and95_i504_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and149_i531_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and115_i520_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and130_i526_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_186to187_bb2_and149_i531_0_stall_in_1_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_cmp37_i471_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2__26_i484_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add192_i548_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_and17_i460_consumed_2_NO_SHIFT_REG <= 1'b0;
		local_bb2_var__u157_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_cmp37_i471_consumed_1_NO_SHIFT_REG <= (local_bb2_add192_i548_inputs_ready & (local_bb2_cmp37_i471_consumed_1_NO_SHIFT_REG | ~(local_bb2_cmp37_i471_stall_in_1)) & local_bb2_add192_i548_stall_local);
		local_bb2__26_i484_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i548_inputs_ready & (local_bb2__26_i484_consumed_0_NO_SHIFT_REG | ~(local_bb2__26_i484_stall_in)) & local_bb2_add192_i548_stall_local);
		local_bb2_add192_i548_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i548_inputs_ready & (local_bb2_add192_i548_consumed_0_NO_SHIFT_REG | ~(local_bb2_add192_i548_stall_in)) & local_bb2_add192_i548_stall_local);
		local_bb2_and17_i460_consumed_2_NO_SHIFT_REG <= (local_bb2_add192_i548_inputs_ready & (local_bb2_and17_i460_consumed_2_NO_SHIFT_REG | ~(local_bb2_and17_i460_stall_in_2)) & local_bb2_add192_i548_stall_local);
		local_bb2_var__u157_consumed_0_NO_SHIFT_REG <= (local_bb2_add192_i548_inputs_ready & (local_bb2_var__u157_consumed_0_NO_SHIFT_REG | ~(local_bb2_var__u157_stall_in)) & local_bb2_add192_i548_stall_local);
	end
end


// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_187to189_bb2_cmp37_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_1_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_2_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_valid_out_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_stall_in_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_187to189_bb2_cmp37_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to189_bb2_cmp37_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to189_bb2_cmp37_i_0_stall_in_0_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_187to189_bb2_cmp37_i_0_valid_out_0_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_187to189_bb2_cmp37_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_cmp37_i),
	.data_out(rnode_187to189_bb2_cmp37_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_187to189_bb2_cmp37_i_0_reg_189_fifo.DEPTH = 2;
defparam rnode_187to189_bb2_cmp37_i_0_reg_189_fifo.DATA_WIDTH = 1;
defparam rnode_187to189_bb2_cmp37_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to189_bb2_cmp37_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_187to189_bb2_cmp37_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp37_i_stall_in_1 = 1'b0;
assign rnode_187to189_bb2_cmp37_i_0_stall_in_0_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_cmp37_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_187to189_bb2_cmp37_i_0_NO_SHIFT_REG = rnode_187to189_bb2_cmp37_i_0_reg_189_NO_SHIFT_REG;
assign rnode_187to189_bb2_cmp37_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_187to189_bb2_cmp37_i_1_NO_SHIFT_REG = rnode_187to189_bb2_cmp37_i_0_reg_189_NO_SHIFT_REG;
assign rnode_187to189_bb2_cmp37_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_187to189_bb2_cmp37_i_2_NO_SHIFT_REG = rnode_187to189_bb2_cmp37_i_0_reg_189_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb2__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb2__26_i_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb2__26_i_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb2__26_i_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb2__26_i_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb2__26_i_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb2__26_i),
	.data_out(rnode_187to188_bb2__26_i_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb2__26_i_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb2__26_i_0_reg_188_fifo.DATA_WIDTH = 1;
defparam rnode_187to188_bb2__26_i_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb2__26_i_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb2__26_i_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__26_i_stall_in = 1'b0;
assign rnode_187to188_bb2__26_i_0_NO_SHIFT_REG = rnode_187to188_bb2__26_i_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2__26_i_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb2__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb2_add192_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i_1_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i_2_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i_3_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_valid_out_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_stall_in_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb2_add192_i_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb2_add192_i_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb2_add192_i_0_stall_in_0_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb2_add192_i_0_valid_out_0_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb2_add192_i_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb2_add192_i),
	.data_out(rnode_187to188_bb2_add192_i_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb2_add192_i_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb2_add192_i_0_reg_188_fifo.DATA_WIDTH = 32;
defparam rnode_187to188_bb2_add192_i_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb2_add192_i_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb2_add192_i_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add192_i_stall_in = 1'b0;
assign rnode_187to188_bb2_add192_i_0_stall_in_0_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb2_add192_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_add192_i_0_NO_SHIFT_REG = rnode_187to188_bb2_add192_i_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_add192_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_add192_i_1_NO_SHIFT_REG = rnode_187to188_bb2_add192_i_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_add192_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_add192_i_2_NO_SHIFT_REG = rnode_187to188_bb2_add192_i_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_add192_i_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_add192_i_3_NO_SHIFT_REG = rnode_187to188_bb2_add192_i_0_reg_188_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_187to189_bb2_and17_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to189_bb2_and17_i_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to189_bb2_and17_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_187to189_bb2_and17_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to189_bb2_and17_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to189_bb2_and17_i_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_187to189_bb2_and17_i_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_187to189_bb2_and17_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_and17_i),
	.data_out(rnode_187to189_bb2_and17_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_187to189_bb2_and17_i_0_reg_189_fifo.DEPTH = 2;
defparam rnode_187to189_bb2_and17_i_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_187to189_bb2_and17_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to189_bb2_and17_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_187to189_bb2_and17_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and17_i_stall_in_2 = 1'b0;
assign rnode_187to189_bb2_and17_i_0_NO_SHIFT_REG = rnode_187to189_bb2_and17_i_0_reg_189_NO_SHIFT_REG;
assign rnode_187to189_bb2_and17_i_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_and17_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb2_var__u156_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u156_0_stall_in_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u156_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u156_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u156_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u156_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u156_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u156_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb2_var__u156_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb2_var__u156_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb2_var__u156_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb2_var__u156_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb2_var__u156_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb2_var__u156),
	.data_out(rnode_187to188_bb2_var__u156_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb2_var__u156_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb2_var__u156_0_reg_188_fifo.DATA_WIDTH = 1;
defparam rnode_187to188_bb2_var__u156_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb2_var__u156_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb2_var__u156_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u156_stall_in = 1'b0;
assign rnode_187to188_bb2_var__u156_0_NO_SHIFT_REG = rnode_187to188_bb2_var__u156_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_var__u156_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb2_var__u156_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_187to189_bb2_cmp37_i471_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_1_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_2_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_valid_out_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_stall_in_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_cmp37_i471_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_187to189_bb2_cmp37_i471_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to189_bb2_cmp37_i471_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to189_bb2_cmp37_i471_0_stall_in_0_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_187to189_bb2_cmp37_i471_0_valid_out_0_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_187to189_bb2_cmp37_i471_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_cmp37_i471),
	.data_out(rnode_187to189_bb2_cmp37_i471_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_187to189_bb2_cmp37_i471_0_reg_189_fifo.DEPTH = 2;
defparam rnode_187to189_bb2_cmp37_i471_0_reg_189_fifo.DATA_WIDTH = 1;
defparam rnode_187to189_bb2_cmp37_i471_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to189_bb2_cmp37_i471_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_187to189_bb2_cmp37_i471_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp37_i471_stall_in_1 = 1'b0;
assign rnode_187to189_bb2_cmp37_i471_0_stall_in_0_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_cmp37_i471_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_187to189_bb2_cmp37_i471_0_NO_SHIFT_REG = rnode_187to189_bb2_cmp37_i471_0_reg_189_NO_SHIFT_REG;
assign rnode_187to189_bb2_cmp37_i471_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_187to189_bb2_cmp37_i471_1_NO_SHIFT_REG = rnode_187to189_bb2_cmp37_i471_0_reg_189_NO_SHIFT_REG;
assign rnode_187to189_bb2_cmp37_i471_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_187to189_bb2_cmp37_i471_2_NO_SHIFT_REG = rnode_187to189_bb2_cmp37_i471_0_reg_189_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb2__26_i484_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i484_0_stall_in_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i484_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i484_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i484_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i484_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i484_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2__26_i484_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb2__26_i484_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb2__26_i484_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb2__26_i484_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb2__26_i484_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb2__26_i484_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb2__26_i484),
	.data_out(rnode_187to188_bb2__26_i484_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb2__26_i484_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb2__26_i484_0_reg_188_fifo.DATA_WIDTH = 1;
defparam rnode_187to188_bb2__26_i484_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb2__26_i484_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb2__26_i484_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__26_i484_stall_in = 1'b0;
assign rnode_187to188_bb2__26_i484_0_NO_SHIFT_REG = rnode_187to188_bb2__26_i484_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2__26_i484_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb2__26_i484_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb2_add192_i548_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i548_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i548_1_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i548_2_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_valid_out_3_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_stall_in_3_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i548_3_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to188_bb2_add192_i548_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_valid_out_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_stall_in_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_add192_i548_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb2_add192_i548_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb2_add192_i548_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb2_add192_i548_0_stall_in_0_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb2_add192_i548_0_valid_out_0_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb2_add192_i548_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb2_add192_i548),
	.data_out(rnode_187to188_bb2_add192_i548_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb2_add192_i548_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb2_add192_i548_0_reg_188_fifo.DATA_WIDTH = 32;
defparam rnode_187to188_bb2_add192_i548_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb2_add192_i548_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb2_add192_i548_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add192_i548_stall_in = 1'b0;
assign rnode_187to188_bb2_add192_i548_0_stall_in_0_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb2_add192_i548_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_add192_i548_0_NO_SHIFT_REG = rnode_187to188_bb2_add192_i548_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_add192_i548_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_add192_i548_1_NO_SHIFT_REG = rnode_187to188_bb2_add192_i548_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_add192_i548_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_add192_i548_2_NO_SHIFT_REG = rnode_187to188_bb2_add192_i548_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_add192_i548_0_valid_out_3_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_add192_i548_3_NO_SHIFT_REG = rnode_187to188_bb2_add192_i548_0_reg_188_NO_SHIFT_REG;

// Register node:
//  * latency = 2
//  * capacity = 2
 logic rnode_187to189_bb2_and17_i460_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i460_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_187to189_bb2_and17_i460_0_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i460_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_187to189_bb2_and17_i460_0_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i460_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i460_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_187to189_bb2_and17_i460_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_187to189_bb2_and17_i460_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to189_bb2_and17_i460_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to189_bb2_and17_i460_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_187to189_bb2_and17_i460_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_187to189_bb2_and17_i460_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_and17_i460),
	.data_out(rnode_187to189_bb2_and17_i460_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_187to189_bb2_and17_i460_0_reg_189_fifo.DEPTH = 2;
defparam rnode_187to189_bb2_and17_i460_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_187to189_bb2_and17_i460_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to189_bb2_and17_i460_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_187to189_bb2_and17_i460_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and17_i460_stall_in_2 = 1'b0;
assign rnode_187to189_bb2_and17_i460_0_NO_SHIFT_REG = rnode_187to189_bb2_and17_i460_0_reg_189_NO_SHIFT_REG;
assign rnode_187to189_bb2_and17_i460_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_and17_i460_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_187to188_bb2_var__u157_0_valid_out_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u157_0_stall_in_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u157_0_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u157_0_reg_188_inputs_ready_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u157_0_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u157_0_valid_out_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u157_0_stall_in_reg_188_NO_SHIFT_REG;
 logic rnode_187to188_bb2_var__u157_0_stall_out_reg_188_NO_SHIFT_REG;

acl_data_fifo rnode_187to188_bb2_var__u157_0_reg_188_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_187to188_bb2_var__u157_0_reg_188_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_187to188_bb2_var__u157_0_stall_in_reg_188_NO_SHIFT_REG),
	.valid_out(rnode_187to188_bb2_var__u157_0_valid_out_reg_188_NO_SHIFT_REG),
	.stall_out(rnode_187to188_bb2_var__u157_0_stall_out_reg_188_NO_SHIFT_REG),
	.data_in(local_bb2_var__u157),
	.data_out(rnode_187to188_bb2_var__u157_0_reg_188_NO_SHIFT_REG)
);

defparam rnode_187to188_bb2_var__u157_0_reg_188_fifo.DEPTH = 1;
defparam rnode_187to188_bb2_var__u157_0_reg_188_fifo.DATA_WIDTH = 1;
defparam rnode_187to188_bb2_var__u157_0_reg_188_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_187to188_bb2_var__u157_0_reg_188_fifo.IMPL = "shift_reg";

assign rnode_187to188_bb2_var__u157_0_reg_188_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u157_stall_in = 1'b0;
assign rnode_187to188_bb2_var__u157_0_NO_SHIFT_REG = rnode_187to188_bb2_var__u157_0_reg_188_NO_SHIFT_REG;
assign rnode_187to188_bb2_var__u157_0_stall_in_reg_188_NO_SHIFT_REG = 1'b0;
assign rnode_187to188_bb2_var__u157_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_not_cmp37_i_stall_local;
wire local_bb2_not_cmp37_i;

assign local_bb2_not_cmp37_i = (rnode_187to189_bb2_cmp37_i_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2__26_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2__26_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2__26_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2__26_i_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2__26_i_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2__26_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(rnode_187to188_bb2__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_188to189_bb2__26_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2__26_i_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2__26_i_0_reg_189_fifo.DATA_WIDTH = 1;
defparam rnode_188to189_bb2__26_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2__26_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2__26_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__26_i_0_NO_SHIFT_REG = rnode_188to189_bb2__26_i_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2__26_i_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__26_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and193_i_valid_out;
wire local_bb2_and193_i_stall_in;
wire local_bb2_and193_i_inputs_ready;
wire local_bb2_and193_i_stall_local;
wire [31:0] local_bb2_and193_i;

assign local_bb2_and193_i_inputs_ready = rnode_187to188_bb2_add192_i_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_and193_i = (rnode_187to188_bb2_add192_i_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb2_and193_i_valid_out = 1'b1;
assign rnode_187to188_bb2_add192_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and195_i_valid_out;
wire local_bb2_and195_i_stall_in;
wire local_bb2_and195_i_inputs_ready;
wire local_bb2_and195_i_stall_local;
wire [31:0] local_bb2_and195_i;

assign local_bb2_and195_i_inputs_ready = rnode_187to188_bb2_add192_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and195_i = (rnode_187to188_bb2_add192_i_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb2_and195_i_valid_out = 1'b1;
assign rnode_187to188_bb2_add192_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and198_i_valid_out;
wire local_bb2_and198_i_stall_in;
wire local_bb2_and198_i_inputs_ready;
wire local_bb2_and198_i_stall_local;
wire [31:0] local_bb2_and198_i;

assign local_bb2_and198_i_inputs_ready = rnode_187to188_bb2_add192_i_0_valid_out_2_NO_SHIFT_REG;
assign local_bb2_and198_i = (rnode_187to188_bb2_add192_i_2_NO_SHIFT_REG & 32'h1);
assign local_bb2_and198_i_valid_out = 1'b1;
assign rnode_187to188_bb2_add192_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and201_i_stall_local;
wire [31:0] local_bb2_and201_i;

assign local_bb2_and201_i = (rnode_187to188_bb2_add192_i_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_var__u156_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u156_0_stall_in_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u156_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u156_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u156_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u156_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u156_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u156_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_var__u156_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_var__u156_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_var__u156_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_var__u156_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_var__u156_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(rnode_187to188_bb2_var__u156_0_NO_SHIFT_REG),
	.data_out(rnode_188to189_bb2_var__u156_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_var__u156_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_var__u156_0_reg_189_fifo.DATA_WIDTH = 1;
defparam rnode_188to189_bb2_var__u156_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_var__u156_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_var__u156_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_var__u156_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_var__u156_0_NO_SHIFT_REG = rnode_188to189_bb2_var__u156_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_var__u156_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_var__u156_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_not_cmp37_i577_stall_local;
wire local_bb2_not_cmp37_i577;

assign local_bb2_not_cmp37_i577 = (rnode_187to189_bb2_cmp37_i471_1_NO_SHIFT_REG ^ 1'b1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2__26_i484_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i484_0_stall_in_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i484_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i484_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i484_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i484_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i484_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__26_i484_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2__26_i484_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2__26_i484_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2__26_i484_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2__26_i484_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2__26_i484_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(rnode_187to188_bb2__26_i484_0_NO_SHIFT_REG),
	.data_out(rnode_188to189_bb2__26_i484_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2__26_i484_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2__26_i484_0_reg_189_fifo.DATA_WIDTH = 1;
defparam rnode_188to189_bb2__26_i484_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2__26_i484_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2__26_i484_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2__26_i484_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__26_i484_0_NO_SHIFT_REG = rnode_188to189_bb2__26_i484_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2__26_i484_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__26_i484_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_and193_i549_valid_out;
wire local_bb2_and193_i549_stall_in;
wire local_bb2_and193_i549_inputs_ready;
wire local_bb2_and193_i549_stall_local;
wire [31:0] local_bb2_and193_i549;

assign local_bb2_and193_i549_inputs_ready = rnode_187to188_bb2_add192_i548_0_valid_out_0_NO_SHIFT_REG;
assign local_bb2_and193_i549 = (rnode_187to188_bb2_add192_i548_0_NO_SHIFT_REG & 32'hFFFFFFF);
assign local_bb2_and193_i549_valid_out = 1'b1;
assign rnode_187to188_bb2_add192_i548_0_stall_in_0_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and195_i550_valid_out;
wire local_bb2_and195_i550_stall_in;
wire local_bb2_and195_i550_inputs_ready;
wire local_bb2_and195_i550_stall_local;
wire [31:0] local_bb2_and195_i550;

assign local_bb2_and195_i550_inputs_ready = rnode_187to188_bb2_add192_i548_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_and195_i550 = (rnode_187to188_bb2_add192_i548_1_NO_SHIFT_REG >> 32'h1B);
assign local_bb2_and195_i550_valid_out = 1'b1;
assign rnode_187to188_bb2_add192_i548_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and198_i551_valid_out;
wire local_bb2_and198_i551_stall_in;
wire local_bb2_and198_i551_inputs_ready;
wire local_bb2_and198_i551_stall_local;
wire [31:0] local_bb2_and198_i551;

assign local_bb2_and198_i551_inputs_ready = rnode_187to188_bb2_add192_i548_0_valid_out_2_NO_SHIFT_REG;
assign local_bb2_and198_i551 = (rnode_187to188_bb2_add192_i548_2_NO_SHIFT_REG & 32'h1);
assign local_bb2_and198_i551_valid_out = 1'b1;
assign rnode_187to188_bb2_add192_i548_0_stall_in_2_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_and201_i552_stall_local;
wire [31:0] local_bb2_and201_i552;

assign local_bb2_and201_i552 = (rnode_187to188_bb2_add192_i548_3_NO_SHIFT_REG & 32'h7FFFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_var__u157_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u157_0_stall_in_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u157_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u157_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u157_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u157_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u157_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_var__u157_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_var__u157_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_var__u157_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_var__u157_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_var__u157_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_var__u157_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(rnode_187to188_bb2_var__u157_0_NO_SHIFT_REG),
	.data_out(rnode_188to189_bb2_var__u157_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_var__u157_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_var__u157_0_reg_189_fifo.DATA_WIDTH = 1;
defparam rnode_188to189_bb2_var__u157_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_var__u157_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_var__u157_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_187to188_bb2_var__u157_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_var__u157_0_NO_SHIFT_REG = rnode_188to189_bb2_var__u157_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_var__u157_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_var__u157_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2__26_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_2_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_valid_out_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_stall_in_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2__26_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2__26_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2__26_i_0_stall_in_0_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2__26_i_0_valid_out_0_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2__26_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(rnode_188to189_bb2__26_i_0_NO_SHIFT_REG),
	.data_out(rnode_189to190_bb2__26_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2__26_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2__26_i_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2__26_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2__26_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2__26_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2__26_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i_0_stall_in_0_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2__26_i_0_NO_SHIFT_REG = rnode_189to190_bb2__26_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2__26_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2__26_i_1_NO_SHIFT_REG = rnode_189to190_bb2__26_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2__26_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2__26_i_2_NO_SHIFT_REG = rnode_189to190_bb2__26_i_0_reg_190_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_and193_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and193_i_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and193_i_1_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and193_i_2_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and193_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_valid_out_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_stall_in_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_and193_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_and193_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_and193_i_0_stall_in_0_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_and193_i_0_valid_out_0_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_and193_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_and193_i),
	.data_out(rnode_188to189_bb2_and193_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_and193_i_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_and193_i_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2_and193_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_and193_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_and193_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and193_i_stall_in = 1'b0;
assign rnode_188to189_bb2_and193_i_0_stall_in_0_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and193_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_and193_i_0_NO_SHIFT_REG = rnode_188to189_bb2_and193_i_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and193_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_and193_i_1_NO_SHIFT_REG = rnode_188to189_bb2_and193_i_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and193_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_and193_i_2_NO_SHIFT_REG = rnode_188to189_bb2_and193_i_0_reg_189_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_and195_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and195_i_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and195_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_and195_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_and195_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_and195_i_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_and195_i_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_and195_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_and195_i),
	.data_out(rnode_188to189_bb2_and195_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_and195_i_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_and195_i_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2_and195_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_and195_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_and195_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and195_i_stall_in = 1'b0;
assign rnode_188to189_bb2_and195_i_0_NO_SHIFT_REG = rnode_188to189_bb2_and195_i_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and195_i_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and195_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_and198_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and198_i_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and198_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_and198_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_and198_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_and198_i_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_and198_i_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_and198_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_and198_i),
	.data_out(rnode_188to189_bb2_and198_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_and198_i_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_and198_i_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2_and198_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_and198_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_and198_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and198_i_stall_in = 1'b0;
assign rnode_188to189_bb2_and198_i_0_NO_SHIFT_REG = rnode_188to189_bb2_and198_i_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and198_i_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and198_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i75_stall_local;
wire [31:0] local_bb2_shr_i_i75;

assign local_bb2_shr_i_i75 = (local_bb2_and201_i >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_var__u156_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u156_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u156_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u156_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u156_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u156_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u156_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u156_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_var__u156_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_var__u156_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_var__u156_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_var__u156_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_var__u156_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(rnode_188to189_bb2_var__u156_0_NO_SHIFT_REG),
	.data_out(rnode_189to190_bb2_var__u156_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_var__u156_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_var__u156_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_var__u156_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_var__u156_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_var__u156_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_var__u156_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_var__u156_0_NO_SHIFT_REG = rnode_189to190_bb2_var__u156_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_var__u156_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_var__u156_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2__26_i484_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_stall_in_2_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_2_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_valid_out_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_stall_in_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__26_i484_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2__26_i484_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2__26_i484_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2__26_i484_0_stall_in_0_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2__26_i484_0_valid_out_0_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2__26_i484_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(rnode_188to189_bb2__26_i484_0_NO_SHIFT_REG),
	.data_out(rnode_189to190_bb2__26_i484_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2__26_i484_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2__26_i484_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2__26_i484_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2__26_i484_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2__26_i484_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2__26_i484_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i484_0_stall_in_0_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i484_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2__26_i484_0_NO_SHIFT_REG = rnode_189to190_bb2__26_i484_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2__26_i484_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2__26_i484_1_NO_SHIFT_REG = rnode_189to190_bb2__26_i484_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2__26_i484_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2__26_i484_2_NO_SHIFT_REG = rnode_189to190_bb2__26_i484_0_reg_190_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_and193_i549_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and193_i549_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and193_i549_1_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and193_i549_2_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and193_i549_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_valid_out_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_stall_in_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and193_i549_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_and193_i549_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_and193_i549_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_and193_i549_0_stall_in_0_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_and193_i549_0_valid_out_0_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_and193_i549_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_and193_i549),
	.data_out(rnode_188to189_bb2_and193_i549_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_and193_i549_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_and193_i549_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2_and193_i549_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_and193_i549_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_and193_i549_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and193_i549_stall_in = 1'b0;
assign rnode_188to189_bb2_and193_i549_0_stall_in_0_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and193_i549_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_and193_i549_0_NO_SHIFT_REG = rnode_188to189_bb2_and193_i549_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and193_i549_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_and193_i549_1_NO_SHIFT_REG = rnode_188to189_bb2_and193_i549_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and193_i549_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_and193_i549_2_NO_SHIFT_REG = rnode_188to189_bb2_and193_i549_0_reg_189_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_and195_i550_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i550_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and195_i550_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i550_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and195_i550_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i550_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i550_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and195_i550_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_and195_i550_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_and195_i550_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_and195_i550_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_and195_i550_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_and195_i550_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_and195_i550),
	.data_out(rnode_188to189_bb2_and195_i550_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_and195_i550_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_and195_i550_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2_and195_i550_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_and195_i550_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_and195_i550_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and195_i550_stall_in = 1'b0;
assign rnode_188to189_bb2_and195_i550_0_NO_SHIFT_REG = rnode_188to189_bb2_and195_i550_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and195_i550_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and195_i550_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2_and198_i551_0_valid_out_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i551_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and198_i551_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i551_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2_and198_i551_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i551_0_valid_out_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i551_0_stall_in_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2_and198_i551_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2_and198_i551_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2_and198_i551_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2_and198_i551_0_stall_in_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2_and198_i551_0_valid_out_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2_and198_i551_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2_and198_i551),
	.data_out(rnode_188to189_bb2_and198_i551_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2_and198_i551_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2_and198_i551_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2_and198_i551_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2_and198_i551_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2_and198_i551_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and198_i551_stall_in = 1'b0;
assign rnode_188to189_bb2_and198_i551_0_NO_SHIFT_REG = rnode_188to189_bb2_and198_i551_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2_and198_i551_0_stall_in_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and198_i551_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_shr_i_i553_stall_local;
wire [31:0] local_bb2_shr_i_i553;

assign local_bb2_shr_i_i553 = (local_bb2_and201_i552 >> 32'h1);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_var__u157_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u157_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u157_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u157_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u157_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u157_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u157_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_var__u157_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_var__u157_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_var__u157_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_var__u157_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_var__u157_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_var__u157_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(rnode_188to189_bb2_var__u157_0_NO_SHIFT_REG),
	.data_out(rnode_189to190_bb2_var__u157_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_var__u157_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_var__u157_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_var__u157_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_var__u157_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_var__u157_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2_var__u157_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_var__u157_0_NO_SHIFT_REG = rnode_189to190_bb2_var__u157_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_var__u157_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_var__u157_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_cond292_i_stall_local;
wire [31:0] local_bb2_cond292_i;

assign local_bb2_cond292_i = (rnode_189to190_bb2__26_i_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u168_stall_local;
wire [31:0] local_bb2_var__u168;

assign local_bb2_var__u168[31:1] = 31'h0;
assign local_bb2_var__u168[0] = rnode_189to190_bb2__26_i_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr216_i_stall_local;
wire [31:0] local_bb2_shr216_i;

assign local_bb2_shr216_i = (rnode_188to189_bb2_and193_i_1_NO_SHIFT_REG >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__pre_i_stall_local;
wire [31:0] local_bb2__pre_i;

assign local_bb2__pre_i = (rnode_188to189_bb2_and195_i_0_NO_SHIFT_REG & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i76_stall_local;
wire [31:0] local_bb2_or_i_i76;

assign local_bb2_or_i_i76 = (local_bb2_shr_i_i75 | local_bb2_and201_i);

// This section implements an unregistered operation.
// 
wire local_bb2_cond292_i611_stall_local;
wire [31:0] local_bb2_cond292_i611;

assign local_bb2_cond292_i611 = (rnode_189to190_bb2__26_i484_1_NO_SHIFT_REG ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u169_stall_local;
wire [31:0] local_bb2_var__u169;

assign local_bb2_var__u169[31:1] = 31'h0;
assign local_bb2_var__u169[0] = rnode_189to190_bb2__26_i484_2_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shr216_i574_stall_local;
wire [31:0] local_bb2_shr216_i574;

assign local_bb2_shr216_i574 = (rnode_188to189_bb2_and193_i549_1_NO_SHIFT_REG >> 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2__pre_i572_stall_local;
wire [31:0] local_bb2__pre_i572;

assign local_bb2__pre_i572 = (rnode_188to189_bb2_and195_i550_0_NO_SHIFT_REG & 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or_i_i554_stall_local;
wire [31:0] local_bb2_or_i_i554;

assign local_bb2_or_i_i554 = (local_bb2_shr_i_i553 | local_bb2_and201_i552);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext_i_stall_local;
wire [31:0] local_bb2_lnot_ext_i;

assign local_bb2_lnot_ext_i = (local_bb2_var__u168 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or219_i_stall_local;
wire [31:0] local_bb2_or219_i;

assign local_bb2_or219_i = (local_bb2_shr216_i | rnode_188to189_bb2_and198_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool213_i_stall_local;
wire local_bb2_tobool213_i;

assign local_bb2_tobool213_i = (local_bb2__pre_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shr1_i_i_stall_local;
wire [31:0] local_bb2_shr1_i_i;

assign local_bb2_shr1_i_i = (local_bb2_or_i_i76 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext_i621_stall_local;
wire [31:0] local_bb2_lnot_ext_i621;

assign local_bb2_lnot_ext_i621 = (local_bb2_var__u169 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or219_i575_stall_local;
wire [31:0] local_bb2_or219_i575;

assign local_bb2_or219_i575 = (local_bb2_shr216_i574 | rnode_188to189_bb2_and198_i551_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_tobool213_i573_stall_local;
wire local_bb2_tobool213_i573;

assign local_bb2_tobool213_i573 = (local_bb2__pre_i572 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_shr1_i_i555_stall_local;
wire [31:0] local_bb2_shr1_i_i555;

assign local_bb2_shr1_i_i555 = (local_bb2_or_i_i554 >> 32'h2);

// This section implements an unregistered operation.
// 
wire local_bb2__40_demorgan_i_stall_local;
wire local_bb2__40_demorgan_i;

assign local_bb2__40_demorgan_i = (rnode_187to189_bb2_cmp37_i_0_NO_SHIFT_REG | local_bb2_tobool213_i);

// This section implements an unregistered operation.
// 
wire local_bb2__42_i_stall_local;
wire local_bb2__42_i;

assign local_bb2__42_i = (local_bb2_tobool213_i & local_bb2_not_cmp37_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or2_i_i_stall_local;
wire [31:0] local_bb2_or2_i_i;

assign local_bb2_or2_i_i = (local_bb2_shr1_i_i | local_bb2_or_i_i76);

// This section implements an unregistered operation.
// 
wire local_bb2__40_demorgan_i576_stall_local;
wire local_bb2__40_demorgan_i576;

assign local_bb2__40_demorgan_i576 = (rnode_187to189_bb2_cmp37_i471_0_NO_SHIFT_REG | local_bb2_tobool213_i573);

// This section implements an unregistered operation.
// 
wire local_bb2__42_i578_stall_local;
wire local_bb2__42_i578;

assign local_bb2__42_i578 = (local_bb2_tobool213_i573 & local_bb2_not_cmp37_i577);

// This section implements an unregistered operation.
// 
wire local_bb2_or2_i_i556_stall_local;
wire [31:0] local_bb2_or2_i_i556;

assign local_bb2_or2_i_i556 = (local_bb2_shr1_i_i555 | local_bb2_or_i_i554);

// This section implements an unregistered operation.
// 
wire local_bb2__43_i_stall_local;
wire [31:0] local_bb2__43_i;

assign local_bb2__43_i = (local_bb2__42_i ? 32'h0 : local_bb2__pre_i);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_i_stall_local;
wire [31:0] local_bb2_shr3_i_i;

assign local_bb2_shr3_i_i = (local_bb2_or2_i_i >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2__43_i579_stall_local;
wire [31:0] local_bb2__43_i579;

assign local_bb2__43_i579 = (local_bb2__42_i578 ? 32'h0 : local_bb2__pre_i572);

// This section implements an unregistered operation.
// 
wire local_bb2_shr3_i_i557_stall_local;
wire [31:0] local_bb2_shr3_i_i557;

assign local_bb2_shr3_i_i557 = (local_bb2_or2_i_i556 >> 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_or4_i_i_stall_local;
wire [31:0] local_bb2_or4_i_i;

assign local_bb2_or4_i_i = (local_bb2_shr3_i_i | local_bb2_or2_i_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or4_i_i558_stall_local;
wire [31:0] local_bb2_or4_i_i558;

assign local_bb2_or4_i_i558 = (local_bb2_shr3_i_i557 | local_bb2_or2_i_i556);

// This section implements an unregistered operation.
// 
wire local_bb2_shr5_i_i_stall_local;
wire [31:0] local_bb2_shr5_i_i;

assign local_bb2_shr5_i_i = (local_bb2_or4_i_i >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_shr5_i_i559_stall_local;
wire [31:0] local_bb2_shr5_i_i559;

assign local_bb2_shr5_i_i559 = (local_bb2_or4_i_i558 >> 32'h8);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_i_i_stall_local;
wire [31:0] local_bb2_or6_i_i;

assign local_bb2_or6_i_i = (local_bb2_shr5_i_i | local_bb2_or4_i_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_i_i560_stall_local;
wire [31:0] local_bb2_or6_i_i560;

assign local_bb2_or6_i_i560 = (local_bb2_shr5_i_i559 | local_bb2_or4_i_i558);

// This section implements an unregistered operation.
// 
wire local_bb2_shr7_i_i_stall_local;
wire [31:0] local_bb2_shr7_i_i;

assign local_bb2_shr7_i_i = (local_bb2_or6_i_i >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_masked_i_i_stall_local;
wire [31:0] local_bb2_or6_masked_i_i;

assign local_bb2_or6_masked_i_i = (local_bb2_or6_i_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_shr7_i_i561_stall_local;
wire [31:0] local_bb2_shr7_i_i561;

assign local_bb2_shr7_i_i561 = (local_bb2_or6_i_i560 >> 32'h10);

// This section implements an unregistered operation.
// 
wire local_bb2_or6_masked_i_i562_stall_local;
wire [31:0] local_bb2_or6_masked_i_i562;

assign local_bb2_or6_masked_i_i562 = (local_bb2_or6_i_i560 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_neg_i_i_stall_local;
wire [31:0] local_bb2_neg_i_i;

assign local_bb2_neg_i_i = (local_bb2_or6_masked_i_i | local_bb2_shr7_i_i);

// This section implements an unregistered operation.
// 
wire local_bb2_neg_i_i563_stall_local;
wire [31:0] local_bb2_neg_i_i563;

assign local_bb2_neg_i_i563 = (local_bb2_or6_masked_i_i562 | local_bb2_shr7_i_i561);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_i_stall_local;
wire [31:0] local_bb2_and_i_i;

assign local_bb2_and_i_i = (local_bb2_neg_i_i ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and_i_i564_stall_local;
wire [31:0] local_bb2_and_i_i564;

assign local_bb2_and_i_i564 = (local_bb2_neg_i_i563 ^ 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2__and_i_i_valid_out;
wire local_bb2__and_i_i_stall_in;
wire local_bb2__and_i_i_inputs_ready;
wire local_bb2__and_i_i_stall_local;
wire [31:0] local_bb2__and_i_i;

thirtysix_six_comp local_bb2__and_i_i_popcnt_instance (
	.data(local_bb2_and_i_i),
	.sum(local_bb2__and_i_i)
);


assign local_bb2__and_i_i_inputs_ready = rnode_187to188_bb2_add192_i_0_valid_out_3_NO_SHIFT_REG;
assign local_bb2__and_i_i_valid_out = 1'b1;
assign rnode_187to188_bb2_add192_i_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2__and_i_i564_valid_out;
wire local_bb2__and_i_i564_stall_in;
wire local_bb2__and_i_i564_inputs_ready;
wire local_bb2__and_i_i564_stall_local;
wire [31:0] local_bb2__and_i_i564;

thirtysix_six_comp local_bb2__and_i_i564_popcnt_instance (
	.data(local_bb2_and_i_i564),
	.sum(local_bb2__and_i_i564)
);


assign local_bb2__and_i_i564_inputs_ready = rnode_187to188_bb2_add192_i548_0_valid_out_3_NO_SHIFT_REG;
assign local_bb2__and_i_i564_valid_out = 1'b1;
assign rnode_187to188_bb2_add192_i548_0_stall_in_3_NO_SHIFT_REG = 1'b0;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2__and_i_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2__and_i_i_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2__and_i_i_1_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2__and_i_i_2_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2__and_i_i_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_valid_out_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_stall_in_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2__and_i_i_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2__and_i_i_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2__and_i_i_0_stall_in_0_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2__and_i_i_0_valid_out_0_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2__and_i_i_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2__and_i_i),
	.data_out(rnode_188to189_bb2__and_i_i_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2__and_i_i_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2__and_i_i_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2__and_i_i_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2__and_i_i_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2__and_i_i_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__and_i_i_stall_in = 1'b0;
assign rnode_188to189_bb2__and_i_i_0_stall_in_0_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__and_i_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2__and_i_i_0_NO_SHIFT_REG = rnode_188to189_bb2__and_i_i_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2__and_i_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2__and_i_i_1_NO_SHIFT_REG = rnode_188to189_bb2__and_i_i_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2__and_i_i_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2__and_i_i_2_NO_SHIFT_REG = rnode_188to189_bb2__and_i_i_0_reg_189_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_188to189_bb2__and_i_i564_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_stall_in_0_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2__and_i_i564_0_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_stall_in_1_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2__and_i_i564_1_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_valid_out_2_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_stall_in_2_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2__and_i_i564_2_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_reg_189_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_188to189_bb2__and_i_i564_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_valid_out_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_stall_in_0_reg_189_NO_SHIFT_REG;
 logic rnode_188to189_bb2__and_i_i564_0_stall_out_reg_189_NO_SHIFT_REG;

acl_data_fifo rnode_188to189_bb2__and_i_i564_0_reg_189_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_188to189_bb2__and_i_i564_0_reg_189_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_188to189_bb2__and_i_i564_0_stall_in_0_reg_189_NO_SHIFT_REG),
	.valid_out(rnode_188to189_bb2__and_i_i564_0_valid_out_0_reg_189_NO_SHIFT_REG),
	.stall_out(rnode_188to189_bb2__and_i_i564_0_stall_out_reg_189_NO_SHIFT_REG),
	.data_in(local_bb2__and_i_i564),
	.data_out(rnode_188to189_bb2__and_i_i564_0_reg_189_NO_SHIFT_REG)
);

defparam rnode_188to189_bb2__and_i_i564_0_reg_189_fifo.DEPTH = 1;
defparam rnode_188to189_bb2__and_i_i564_0_reg_189_fifo.DATA_WIDTH = 32;
defparam rnode_188to189_bb2__and_i_i564_0_reg_189_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_188to189_bb2__and_i_i564_0_reg_189_fifo.IMPL = "shift_reg";

assign rnode_188to189_bb2__and_i_i564_0_reg_189_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__and_i_i564_stall_in = 1'b0;
assign rnode_188to189_bb2__and_i_i564_0_stall_in_0_reg_189_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__and_i_i564_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2__and_i_i564_0_NO_SHIFT_REG = rnode_188to189_bb2__and_i_i564_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2__and_i_i564_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2__and_i_i564_1_NO_SHIFT_REG = rnode_188to189_bb2__and_i_i564_0_reg_189_NO_SHIFT_REG;
assign rnode_188to189_bb2__and_i_i564_0_valid_out_2_NO_SHIFT_REG = 1'b1;
assign rnode_188to189_bb2__and_i_i564_2_NO_SHIFT_REG = rnode_188to189_bb2__and_i_i564_0_reg_189_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_and9_i_i_stall_local;
wire [31:0] local_bb2_and9_i_i;

assign local_bb2_and9_i_i = (rnode_188to189_bb2__and_i_i_0_NO_SHIFT_REG & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and203_i_stall_local;
wire [31:0] local_bb2_and203_i;

assign local_bb2_and203_i = (rnode_188to189_bb2__and_i_i_1_NO_SHIFT_REG & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_and206_i_stall_local;
wire [31:0] local_bb2_and206_i;

assign local_bb2_and206_i = (rnode_188to189_bb2__and_i_i_2_NO_SHIFT_REG & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_and9_i_i565_stall_local;
wire [31:0] local_bb2_and9_i_i565;

assign local_bb2_and9_i_i565 = (rnode_188to189_bb2__and_i_i564_0_NO_SHIFT_REG & 32'h1F);

// This section implements an unregistered operation.
// 
wire local_bb2_and203_i566_stall_local;
wire [31:0] local_bb2_and203_i566;

assign local_bb2_and203_i566 = (rnode_188to189_bb2__and_i_i564_1_NO_SHIFT_REG & 32'h18);

// This section implements an unregistered operation.
// 
wire local_bb2_and206_i568_stall_local;
wire [31:0] local_bb2_and206_i568;

assign local_bb2_and206_i568 = (rnode_188to189_bb2__and_i_i564_2_NO_SHIFT_REG & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_sub239_i_stall_local;
wire [31:0] local_bb2_sub239_i;

assign local_bb2_sub239_i = (32'h0 - local_bb2_and9_i_i);

// This section implements an unregistered operation.
// 
wire local_bb2_shl204_i_stall_local;
wire [31:0] local_bb2_shl204_i;

assign local_bb2_shl204_i = (rnode_188to189_bb2_and193_i_0_NO_SHIFT_REG << local_bb2_and203_i);

// This section implements an unregistered operation.
// 
wire local_bb2_sub239_i587_stall_local;
wire [31:0] local_bb2_sub239_i587;

assign local_bb2_sub239_i587 = (32'h0 - local_bb2_and9_i_i565);

// This section implements an unregistered operation.
// 
wire local_bb2_shl204_i567_stall_local;
wire [31:0] local_bb2_shl204_i567;

assign local_bb2_shl204_i567 = (rnode_188to189_bb2_and193_i549_0_NO_SHIFT_REG << local_bb2_and203_i566);

// This section implements an unregistered operation.
// 
wire local_bb2_cond244_i_stall_local;
wire [31:0] local_bb2_cond244_i;

assign local_bb2_cond244_i = (rnode_187to189_bb2_cmp37_i_2_NO_SHIFT_REG ? local_bb2_sub239_i : local_bb2__43_i);

// This section implements an unregistered operation.
// 
wire local_bb2_and205_i_stall_local;
wire [31:0] local_bb2_and205_i;

assign local_bb2_and205_i = (local_bb2_shl204_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond244_i588_stall_local;
wire [31:0] local_bb2_cond244_i588;

assign local_bb2_cond244_i588 = (rnode_187to189_bb2_cmp37_i471_2_NO_SHIFT_REG ? local_bb2_sub239_i587 : local_bb2__43_i579);

// This section implements an unregistered operation.
// 
wire local_bb2_and205_i569_stall_local;
wire [31:0] local_bb2_and205_i569;

assign local_bb2_and205_i569 = (local_bb2_shl204_i567 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_add245_i_stall_local;
wire [31:0] local_bb2_add245_i;

assign local_bb2_add245_i = (local_bb2_cond244_i + rnode_187to189_bb2_and17_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_fold_i77_stall_local;
wire [31:0] local_bb2_fold_i77;

assign local_bb2_fold_i77 = (local_bb2_cond244_i + rnode_187to189_bb2_shr16_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl207_i_stall_local;
wire [31:0] local_bb2_shl207_i;

assign local_bb2_shl207_i = (local_bb2_and205_i << local_bb2_and206_i);

// This section implements an unregistered operation.
// 
wire local_bb2_add245_i589_stall_local;
wire [31:0] local_bb2_add245_i589;

assign local_bb2_add245_i589 = (local_bb2_cond244_i588 + rnode_187to189_bb2_and17_i460_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_fold_i591_stall_local;
wire [31:0] local_bb2_fold_i591;

assign local_bb2_fold_i591 = (local_bb2_cond244_i588 + rnode_187to189_bb2_shr16_i459_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_shl207_i570_stall_local;
wire [31:0] local_bb2_shl207_i570;

assign local_bb2_shl207_i570 = (local_bb2_and205_i569 << local_bb2_and206_i568);

// This section implements an unregistered operation.
// 
wire local_bb2_and247_i_stall_local;
wire [31:0] local_bb2_and247_i;

assign local_bb2_and247_i = (local_bb2_add245_i & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb2_and250_i_stall_local;
wire [31:0] local_bb2_and250_i;

assign local_bb2_and250_i = (local_bb2_fold_i77 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i_stall_local;
wire [31:0] local_bb2_and269_i;

assign local_bb2_and269_i = (local_bb2_fold_i77 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and208_i_stall_local;
wire [31:0] local_bb2_and208_i;

assign local_bb2_and208_i = (local_bb2_shl207_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and247_i590_stall_local;
wire [31:0] local_bb2_and247_i590;

assign local_bb2_and247_i590 = (local_bb2_add245_i589 & 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb2_and250_i592_stall_local;
wire [31:0] local_bb2_and250_i592;

assign local_bb2_and250_i592 = (local_bb2_fold_i591 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i603_stall_local;
wire [31:0] local_bb2_and269_i603;

assign local_bb2_and269_i603 = (local_bb2_fold_i591 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb2_and208_i571_stall_local;
wire [31:0] local_bb2_and208_i571;

assign local_bb2_and208_i571 = (local_bb2_shl207_i570 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_notlhs_i_stall_local;
wire local_bb2_notlhs_i;

assign local_bb2_notlhs_i = (local_bb2_and247_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_notrhs_i_stall_local;
wire local_bb2_notrhs_i;

assign local_bb2_notrhs_i = (local_bb2_and250_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__44_i_stall_local;
wire [31:0] local_bb2__44_i;

assign local_bb2__44_i = (local_bb2__40_demorgan_i ? local_bb2_and208_i : local_bb2_or219_i);

// This section implements an unregistered operation.
// 
wire local_bb2_notlhs_i593_stall_local;
wire local_bb2_notlhs_i593;

assign local_bb2_notlhs_i593 = (local_bb2_and247_i590 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_notrhs_i594_stall_local;
wire local_bb2_notrhs_i594;

assign local_bb2_notrhs_i594 = (local_bb2_and250_i592 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2__44_i580_stall_local;
wire [31:0] local_bb2__44_i580;

assign local_bb2__44_i580 = (local_bb2__40_demorgan_i576 ? local_bb2_and208_i571 : local_bb2_or219_i575);

// This section implements an unregistered operation.
// 
wire local_bb2_not__46_i_stall_local;
wire local_bb2_not__46_i;

assign local_bb2_not__46_i = (local_bb2_notrhs_i | local_bb2_notlhs_i);

// This section implements an unregistered operation.
// 
wire local_bb2__45_i_stall_local;
wire [31:0] local_bb2__45_i;

assign local_bb2__45_i = (local_bb2__42_i ? rnode_188to189_bb2_and193_i_2_NO_SHIFT_REG : local_bb2__44_i);

// This section implements an unregistered operation.
// 
wire local_bb2_not__46_i595_stall_local;
wire local_bb2_not__46_i595;

assign local_bb2_not__46_i595 = (local_bb2_notrhs_i594 | local_bb2_notlhs_i593);

// This section implements an unregistered operation.
// 
wire local_bb2__45_i581_stall_local;
wire [31:0] local_bb2__45_i581;

assign local_bb2__45_i581 = (local_bb2__42_i578 ? rnode_188to189_bb2_and193_i549_2_NO_SHIFT_REG : local_bb2__44_i580);

// This section implements an unregistered operation.
// 
wire local_bb2_and225_i_stall_local;
wire [31:0] local_bb2_and225_i;

assign local_bb2_and225_i = (local_bb2__45_i & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i_stall_local;
wire [31:0] local_bb2_and270_i;

assign local_bb2_and270_i = (local_bb2__45_i & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_shr271_i_stall_local;
wire [31:0] local_bb2_shr271_i;

assign local_bb2_shr271_i = (local_bb2__45_i >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_and225_i582_stall_local;
wire [31:0] local_bb2_and225_i582;

assign local_bb2_and225_i582 = (local_bb2__45_i581 & 32'h7FFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_and270_i600_stall_local;
wire [31:0] local_bb2_and270_i600;

assign local_bb2_and270_i600 = (local_bb2__45_i581 & 32'h7);

// This section implements an unregistered operation.
// 
wire local_bb2_shr271_i601_stall_local;
wire [31:0] local_bb2_shr271_i601;

assign local_bb2_shr271_i601 = (local_bb2__45_i581 >> 32'h3);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_i_stall_local;
wire local_bb2_cmp226_i;

assign local_bb2_cmp226_i = (local_bb2_and225_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp296_i_stall_local;
wire local_bb2_cmp296_i;

assign local_bb2_cmp296_i = (local_bb2_and270_i > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp299_i_stall_local;
wire local_bb2_cmp299_i;

assign local_bb2_cmp299_i = (local_bb2_and270_i == 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_i583_stall_local;
wire local_bb2_cmp226_i583;

assign local_bb2_cmp226_i583 = (local_bb2_and225_i582 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp296_i615_stall_local;
wire local_bb2_cmp296_i615;

assign local_bb2_cmp296_i615 = (local_bb2_and270_i600 > 32'h4);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i603_valid_out;
wire local_bb2_and269_i603_stall_in;
 reg local_bb2_and269_i603_consumed_0_NO_SHIFT_REG;
wire local_bb2_add245_i589_valid_out_1;
wire local_bb2_add245_i589_stall_in_1;
 reg local_bb2_add245_i589_consumed_1_NO_SHIFT_REG;
wire local_bb2_not__46_i595_valid_out;
wire local_bb2_not__46_i595_stall_in;
 reg local_bb2_not__46_i595_consumed_0_NO_SHIFT_REG;
wire local_bb2_not_cmp37_i577_valid_out_1;
wire local_bb2_not_cmp37_i577_stall_in_1;
 reg local_bb2_not_cmp37_i577_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr271_i601_valid_out;
wire local_bb2_shr271_i601_stall_in;
 reg local_bb2_shr271_i601_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp226_i583_valid_out;
wire local_bb2_cmp226_i583_stall_in;
 reg local_bb2_cmp226_i583_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp296_i615_valid_out;
wire local_bb2_cmp296_i615_stall_in;
 reg local_bb2_cmp296_i615_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i616_valid_out;
wire local_bb2_cmp299_i616_stall_in;
 reg local_bb2_cmp299_i616_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i616_inputs_ready;
wire local_bb2_cmp299_i616_stall_local;
wire local_bb2_cmp299_i616;

assign local_bb2_cmp299_i616_inputs_ready = (rnode_187to189_bb2_shr16_i459_0_valid_out_NO_SHIFT_REG & rnode_187to189_bb2_cmp37_i471_0_valid_out_2_NO_SHIFT_REG & rnode_187to189_bb2_and17_i460_0_valid_out_NO_SHIFT_REG & rnode_187to189_bb2_cmp37_i471_0_valid_out_0_NO_SHIFT_REG & rnode_188to189_bb2_and193_i549_0_valid_out_2_NO_SHIFT_REG & rnode_187to189_bb2_cmp37_i471_0_valid_out_1_NO_SHIFT_REG & rnode_188to189_bb2_and195_i550_0_valid_out_NO_SHIFT_REG & rnode_188to189_bb2_and193_i549_0_valid_out_1_NO_SHIFT_REG & rnode_188to189_bb2_and198_i551_0_valid_out_NO_SHIFT_REG & rnode_188to189_bb2_and193_i549_0_valid_out_0_NO_SHIFT_REG & rnode_188to189_bb2__and_i_i564_0_valid_out_1_NO_SHIFT_REG & rnode_188to189_bb2__and_i_i564_0_valid_out_2_NO_SHIFT_REG & rnode_188to189_bb2__and_i_i564_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2_cmp299_i616 = (local_bb2_and270_i600 == 32'h4);
assign local_bb2_and269_i603_valid_out = 1'b1;
assign local_bb2_add245_i589_valid_out_1 = 1'b1;
assign local_bb2_not__46_i595_valid_out = 1'b1;
assign local_bb2_not_cmp37_i577_valid_out_1 = 1'b1;
assign local_bb2_shr271_i601_valid_out = 1'b1;
assign local_bb2_cmp226_i583_valid_out = 1'b1;
assign local_bb2_cmp296_i615_valid_out = 1'b1;
assign local_bb2_cmp299_i616_valid_out = 1'b1;
assign rnode_187to189_bb2_shr16_i459_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_cmp37_i471_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_and17_i460_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_cmp37_i471_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and193_i549_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_cmp37_i471_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and195_i550_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and193_i549_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and198_i551_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and193_i549_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__and_i_i564_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__and_i_i564_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__and_i_i564_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_and269_i603_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add245_i589_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_not__46_i595_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_not_cmp37_i577_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr271_i601_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp226_i583_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp296_i615_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp299_i616_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_and269_i603_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i616_inputs_ready & (local_bb2_and269_i603_consumed_0_NO_SHIFT_REG | ~(local_bb2_and269_i603_stall_in)) & local_bb2_cmp299_i616_stall_local);
		local_bb2_add245_i589_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp299_i616_inputs_ready & (local_bb2_add245_i589_consumed_1_NO_SHIFT_REG | ~(local_bb2_add245_i589_stall_in_1)) & local_bb2_cmp299_i616_stall_local);
		local_bb2_not__46_i595_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i616_inputs_ready & (local_bb2_not__46_i595_consumed_0_NO_SHIFT_REG | ~(local_bb2_not__46_i595_stall_in)) & local_bb2_cmp299_i616_stall_local);
		local_bb2_not_cmp37_i577_consumed_1_NO_SHIFT_REG <= (local_bb2_cmp299_i616_inputs_ready & (local_bb2_not_cmp37_i577_consumed_1_NO_SHIFT_REG | ~(local_bb2_not_cmp37_i577_stall_in_1)) & local_bb2_cmp299_i616_stall_local);
		local_bb2_shr271_i601_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i616_inputs_ready & (local_bb2_shr271_i601_consumed_0_NO_SHIFT_REG | ~(local_bb2_shr271_i601_stall_in)) & local_bb2_cmp299_i616_stall_local);
		local_bb2_cmp226_i583_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i616_inputs_ready & (local_bb2_cmp226_i583_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp226_i583_stall_in)) & local_bb2_cmp299_i616_stall_local);
		local_bb2_cmp296_i615_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i616_inputs_ready & (local_bb2_cmp296_i615_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp296_i615_stall_in)) & local_bb2_cmp299_i616_stall_local);
		local_bb2_cmp299_i616_consumed_0_NO_SHIFT_REG <= (local_bb2_cmp299_i616_inputs_ready & (local_bb2_cmp299_i616_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp299_i616_stall_in)) & local_bb2_cmp299_i616_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_not_i_stall_local;
wire local_bb2_cmp226_not_i;

assign local_bb2_cmp226_not_i = (local_bb2_cmp226_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2_and269_i_valid_out;
wire local_bb2_and269_i_stall_in;
 reg local_bb2_and269_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_add245_i_valid_out_1;
wire local_bb2_add245_i_stall_in_1;
 reg local_bb2_add245_i_consumed_1_NO_SHIFT_REG;
wire local_bb2_not_cmp37_i_valid_out_1;
wire local_bb2_not_cmp37_i_stall_in_1;
 reg local_bb2_not_cmp37_i_consumed_1_NO_SHIFT_REG;
wire local_bb2_shr271_i_valid_out;
wire local_bb2_shr271_i_stall_in;
 reg local_bb2_shr271_i_consumed_0_NO_SHIFT_REG;
wire local_bb2__47_i_valid_out;
wire local_bb2__47_i_stall_in;
 reg local_bb2__47_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp296_i_valid_out;
wire local_bb2_cmp296_i_stall_in;
 reg local_bb2_cmp296_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp299_i_valid_out;
wire local_bb2_cmp299_i_stall_in;
 reg local_bb2_cmp299_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_cmp226_not_i_valid_out;
wire local_bb2_cmp226_not_i_stall_in;
 reg local_bb2_cmp226_not_i_consumed_0_NO_SHIFT_REG;
wire local_bb2__47_i_inputs_ready;
wire local_bb2__47_i_stall_local;
wire local_bb2__47_i;

assign local_bb2__47_i_inputs_ready = (rnode_187to189_bb2_shr16_i_0_valid_out_NO_SHIFT_REG & rnode_187to189_bb2_cmp37_i_0_valid_out_2_NO_SHIFT_REG & rnode_187to189_bb2_and17_i_0_valid_out_NO_SHIFT_REG & rnode_187to189_bb2_cmp37_i_0_valid_out_0_NO_SHIFT_REG & rnode_188to189_bb2_and193_i_0_valid_out_2_NO_SHIFT_REG & rnode_187to189_bb2_cmp37_i_0_valid_out_1_NO_SHIFT_REG & rnode_188to189_bb2_and195_i_0_valid_out_NO_SHIFT_REG & rnode_188to189_bb2_and193_i_0_valid_out_1_NO_SHIFT_REG & rnode_188to189_bb2_and198_i_0_valid_out_NO_SHIFT_REG & rnode_188to189_bb2_and193_i_0_valid_out_0_NO_SHIFT_REG & rnode_188to189_bb2__and_i_i_0_valid_out_1_NO_SHIFT_REG & rnode_188to189_bb2__and_i_i_0_valid_out_2_NO_SHIFT_REG & rnode_188to189_bb2__and_i_i_0_valid_out_0_NO_SHIFT_REG);
assign local_bb2__47_i = (local_bb2_cmp226_i | local_bb2_not__46_i);
assign local_bb2_and269_i_valid_out = 1'b1;
assign local_bb2_add245_i_valid_out_1 = 1'b1;
assign local_bb2_not_cmp37_i_valid_out_1 = 1'b1;
assign local_bb2_shr271_i_valid_out = 1'b1;
assign local_bb2__47_i_valid_out = 1'b1;
assign local_bb2_cmp296_i_valid_out = 1'b1;
assign local_bb2_cmp299_i_valid_out = 1'b1;
assign local_bb2_cmp226_not_i_valid_out = 1'b1;
assign rnode_187to189_bb2_shr16_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_cmp37_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_and17_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_cmp37_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and193_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_187to189_bb2_cmp37_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and195_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and193_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and198_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2_and193_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__and_i_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__and_i_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_188to189_bb2__and_i_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_and269_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_add245_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_not_cmp37_i_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_shr271_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__47_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp296_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp299_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_cmp226_not_i_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_and269_i_consumed_0_NO_SHIFT_REG <= (local_bb2__47_i_inputs_ready & (local_bb2_and269_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_and269_i_stall_in)) & local_bb2__47_i_stall_local);
		local_bb2_add245_i_consumed_1_NO_SHIFT_REG <= (local_bb2__47_i_inputs_ready & (local_bb2_add245_i_consumed_1_NO_SHIFT_REG | ~(local_bb2_add245_i_stall_in_1)) & local_bb2__47_i_stall_local);
		local_bb2_not_cmp37_i_consumed_1_NO_SHIFT_REG <= (local_bb2__47_i_inputs_ready & (local_bb2_not_cmp37_i_consumed_1_NO_SHIFT_REG | ~(local_bb2_not_cmp37_i_stall_in_1)) & local_bb2__47_i_stall_local);
		local_bb2_shr271_i_consumed_0_NO_SHIFT_REG <= (local_bb2__47_i_inputs_ready & (local_bb2_shr271_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_shr271_i_stall_in)) & local_bb2__47_i_stall_local);
		local_bb2__47_i_consumed_0_NO_SHIFT_REG <= (local_bb2__47_i_inputs_ready & (local_bb2__47_i_consumed_0_NO_SHIFT_REG | ~(local_bb2__47_i_stall_in)) & local_bb2__47_i_stall_local);
		local_bb2_cmp296_i_consumed_0_NO_SHIFT_REG <= (local_bb2__47_i_inputs_ready & (local_bb2_cmp296_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp296_i_stall_in)) & local_bb2__47_i_stall_local);
		local_bb2_cmp299_i_consumed_0_NO_SHIFT_REG <= (local_bb2__47_i_inputs_ready & (local_bb2_cmp299_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp299_i_stall_in)) & local_bb2__47_i_stall_local);
		local_bb2_cmp226_not_i_consumed_0_NO_SHIFT_REG <= (local_bb2__47_i_inputs_ready & (local_bb2_cmp226_not_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_cmp226_not_i_stall_in)) & local_bb2__47_i_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_and269_i603_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i603_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_and269_i603_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i603_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_and269_i603_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i603_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i603_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i603_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_and269_i603_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_and269_i603_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_and269_i603_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_and269_i603_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_and269_i603_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_and269_i603),
	.data_out(rnode_189to190_bb2_and269_i603_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_and269_i603_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_and269_i603_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_189to190_bb2_and269_i603_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_and269_i603_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_and269_i603_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and269_i603_stall_in = 1'b0;
assign rnode_189to190_bb2_and269_i603_0_NO_SHIFT_REG = rnode_189to190_bb2_and269_i603_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_and269_i603_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_and269_i603_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_add245_i589_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i589_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_add245_i589_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i589_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_add245_i589_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i589_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i589_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i589_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_add245_i589_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_add245_i589_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_add245_i589_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_add245_i589_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_add245_i589_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_add245_i589),
	.data_out(rnode_189to190_bb2_add245_i589_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_add245_i589_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_add245_i589_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_189to190_bb2_add245_i589_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_add245_i589_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_add245_i589_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add245_i589_stall_in_1 = 1'b0;
assign rnode_189to190_bb2_add245_i589_0_NO_SHIFT_REG = rnode_189to190_bb2_add245_i589_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_add245_i589_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_add245_i589_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_not__46_i595_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not__46_i595_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not__46_i595_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not__46_i595_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not__46_i595_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not__46_i595_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not__46_i595_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not__46_i595_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_not__46_i595_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_not__46_i595_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_not__46_i595_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_not__46_i595_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_not__46_i595_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_not__46_i595),
	.data_out(rnode_189to190_bb2_not__46_i595_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_not__46_i595_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_not__46_i595_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_not__46_i595_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_not__46_i595_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_not__46_i595_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not__46_i595_stall_in = 1'b0;
assign rnode_189to190_bb2_not__46_i595_0_NO_SHIFT_REG = rnode_189to190_bb2_not__46_i595_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_not__46_i595_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_not__46_i595_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_not_cmp37_i577_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i577_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i577_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i577_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i577_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i577_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i577_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i577_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_not_cmp37_i577_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_not_cmp37_i577_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_not_cmp37_i577_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_not_cmp37_i577_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_not_cmp37_i577_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_not_cmp37_i577),
	.data_out(rnode_189to190_bb2_not_cmp37_i577_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_not_cmp37_i577_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_not_cmp37_i577_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_not_cmp37_i577_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_not_cmp37_i577_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_not_cmp37_i577_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not_cmp37_i577_stall_in_1 = 1'b0;
assign rnode_189to190_bb2_not_cmp37_i577_0_NO_SHIFT_REG = rnode_189to190_bb2_not_cmp37_i577_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_not_cmp37_i577_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_not_cmp37_i577_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_shr271_i601_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i601_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_shr271_i601_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i601_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_shr271_i601_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i601_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i601_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i601_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_shr271_i601_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_shr271_i601_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_shr271_i601_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_shr271_i601_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_shr271_i601_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_shr271_i601),
	.data_out(rnode_189to190_bb2_shr271_i601_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_shr271_i601_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_shr271_i601_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_189to190_bb2_shr271_i601_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_shr271_i601_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_shr271_i601_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr271_i601_stall_in = 1'b0;
assign rnode_189to190_bb2_shr271_i601_0_NO_SHIFT_REG = rnode_189to190_bb2_shr271_i601_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_shr271_i601_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_shr271_i601_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_cmp226_i583_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_valid_out_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_stall_in_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_i583_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_cmp226_i583_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_cmp226_i583_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_cmp226_i583_0_stall_in_0_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_cmp226_i583_0_valid_out_0_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_cmp226_i583_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_cmp226_i583),
	.data_out(rnode_189to190_bb2_cmp226_i583_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_cmp226_i583_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_cmp226_i583_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_cmp226_i583_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_cmp226_i583_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_cmp226_i583_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp226_i583_stall_in = 1'b0;
assign rnode_189to190_bb2_cmp226_i583_0_stall_in_0_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp226_i583_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2_cmp226_i583_0_NO_SHIFT_REG = rnode_189to190_bb2_cmp226_i583_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_cmp226_i583_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2_cmp226_i583_1_NO_SHIFT_REG = rnode_189to190_bb2_cmp226_i583_0_reg_190_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_cmp296_i615_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i615_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i615_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i615_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i615_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i615_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i615_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i615_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_cmp296_i615_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_cmp296_i615_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_cmp296_i615_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_cmp296_i615_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_cmp296_i615_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_cmp296_i615),
	.data_out(rnode_189to190_bb2_cmp296_i615_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_cmp296_i615_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_cmp296_i615_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_cmp296_i615_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_cmp296_i615_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_cmp296_i615_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp296_i615_stall_in = 1'b0;
assign rnode_189to190_bb2_cmp296_i615_0_NO_SHIFT_REG = rnode_189to190_bb2_cmp296_i615_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_cmp296_i615_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp296_i615_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_cmp299_i616_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i616_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i616_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i616_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i616_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i616_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i616_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i616_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_cmp299_i616_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_cmp299_i616_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_cmp299_i616_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_cmp299_i616_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_cmp299_i616_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_cmp299_i616),
	.data_out(rnode_189to190_bb2_cmp299_i616_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_cmp299_i616_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_cmp299_i616_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_cmp299_i616_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_cmp299_i616_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_cmp299_i616_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp299_i616_stall_in = 1'b0;
assign rnode_189to190_bb2_cmp299_i616_0_NO_SHIFT_REG = rnode_189to190_bb2_cmp299_i616_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_cmp299_i616_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp299_i616_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_and269_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_and269_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_and269_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_and269_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_and269_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_and269_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_and269_i_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_and269_i_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_and269_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_and269_i),
	.data_out(rnode_189to190_bb2_and269_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_and269_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_and269_i_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_189to190_bb2_and269_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_and269_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_and269_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_and269_i_stall_in = 1'b0;
assign rnode_189to190_bb2_and269_i_0_NO_SHIFT_REG = rnode_189to190_bb2_and269_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_and269_i_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_and269_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_add245_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_add245_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_add245_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_add245_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_add245_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_add245_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_add245_i_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_add245_i_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_add245_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_add245_i),
	.data_out(rnode_189to190_bb2_add245_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_add245_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_add245_i_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_189to190_bb2_add245_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_add245_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_add245_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_add245_i_stall_in_1 = 1'b0;
assign rnode_189to190_bb2_add245_i_0_NO_SHIFT_REG = rnode_189to190_bb2_add245_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_add245_i_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_add245_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_not_cmp37_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_not_cmp37_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_not_cmp37_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_not_cmp37_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_not_cmp37_i_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_not_cmp37_i_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_not_cmp37_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_not_cmp37_i),
	.data_out(rnode_189to190_bb2_not_cmp37_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_not_cmp37_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_not_cmp37_i_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_not_cmp37_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_not_cmp37_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_not_cmp37_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_not_cmp37_i_stall_in_1 = 1'b0;
assign rnode_189to190_bb2_not_cmp37_i_0_NO_SHIFT_REG = rnode_189to190_bb2_not_cmp37_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_not_cmp37_i_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_not_cmp37_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_shr271_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_shr271_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_189to190_bb2_shr271_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_shr271_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_shr271_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_shr271_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_shr271_i_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_shr271_i_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_shr271_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_shr271_i),
	.data_out(rnode_189to190_bb2_shr271_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_shr271_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_shr271_i_0_reg_190_fifo.DATA_WIDTH = 32;
defparam rnode_189to190_bb2_shr271_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_shr271_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_shr271_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_shr271_i_stall_in = 1'b0;
assign rnode_189to190_bb2_shr271_i_0_NO_SHIFT_REG = rnode_189to190_bb2_shr271_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_shr271_i_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_shr271_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2__47_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_valid_out_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_stall_in_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2__47_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2__47_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2__47_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2__47_i_0_stall_in_0_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2__47_i_0_valid_out_0_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2__47_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2__47_i),
	.data_out(rnode_189to190_bb2__47_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2__47_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2__47_i_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2__47_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2__47_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2__47_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__47_i_stall_in = 1'b0;
assign rnode_189to190_bb2__47_i_0_stall_in_0_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__47_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2__47_i_0_NO_SHIFT_REG = rnode_189to190_bb2__47_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2__47_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2__47_i_1_NO_SHIFT_REG = rnode_189to190_bb2__47_i_0_reg_190_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_cmp296_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp296_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_cmp296_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_cmp296_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_cmp296_i_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_cmp296_i_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_cmp296_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_cmp296_i),
	.data_out(rnode_189to190_bb2_cmp296_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_cmp296_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_cmp296_i_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_cmp296_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_cmp296_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_cmp296_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp296_i_stall_in = 1'b0;
assign rnode_189to190_bb2_cmp296_i_0_NO_SHIFT_REG = rnode_189to190_bb2_cmp296_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_cmp296_i_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp296_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_cmp299_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i_0_stall_in_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i_0_valid_out_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i_0_stall_in_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp299_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_cmp299_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_cmp299_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_cmp299_i_0_stall_in_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_cmp299_i_0_valid_out_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_cmp299_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_cmp299_i),
	.data_out(rnode_189to190_bb2_cmp299_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_cmp299_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_cmp299_i_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_cmp299_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_cmp299_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_cmp299_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp299_i_stall_in = 1'b0;
assign rnode_189to190_bb2_cmp299_i_0_NO_SHIFT_REG = rnode_189to190_bb2_cmp299_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_cmp299_i_0_stall_in_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp299_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_189to190_bb2_cmp226_not_i_0_valid_out_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_stall_in_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_valid_out_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_stall_in_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_1_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_reg_190_inputs_ready_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_valid_out_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_stall_in_0_reg_190_NO_SHIFT_REG;
 logic rnode_189to190_bb2_cmp226_not_i_0_stall_out_reg_190_NO_SHIFT_REG;

acl_data_fifo rnode_189to190_bb2_cmp226_not_i_0_reg_190_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_189to190_bb2_cmp226_not_i_0_reg_190_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_189to190_bb2_cmp226_not_i_0_stall_in_0_reg_190_NO_SHIFT_REG),
	.valid_out(rnode_189to190_bb2_cmp226_not_i_0_valid_out_0_reg_190_NO_SHIFT_REG),
	.stall_out(rnode_189to190_bb2_cmp226_not_i_0_stall_out_reg_190_NO_SHIFT_REG),
	.data_in(local_bb2_cmp226_not_i),
	.data_out(rnode_189to190_bb2_cmp226_not_i_0_reg_190_NO_SHIFT_REG)
);

defparam rnode_189to190_bb2_cmp226_not_i_0_reg_190_fifo.DEPTH = 1;
defparam rnode_189to190_bb2_cmp226_not_i_0_reg_190_fifo.DATA_WIDTH = 1;
defparam rnode_189to190_bb2_cmp226_not_i_0_reg_190_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_189to190_bb2_cmp226_not_i_0_reg_190_fifo.IMPL = "shift_reg";

assign rnode_189to190_bb2_cmp226_not_i_0_reg_190_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_cmp226_not_i_stall_in = 1'b0;
assign rnode_189to190_bb2_cmp226_not_i_0_stall_in_0_reg_190_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp226_not_i_0_valid_out_0_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2_cmp226_not_i_0_NO_SHIFT_REG = rnode_189to190_bb2_cmp226_not_i_0_reg_190_NO_SHIFT_REG;
assign rnode_189to190_bb2_cmp226_not_i_0_valid_out_1_NO_SHIFT_REG = 1'b1;
assign rnode_189to190_bb2_cmp226_not_i_1_NO_SHIFT_REG = rnode_189to190_bb2_cmp226_not_i_0_reg_190_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shl273_i604_stall_local;
wire [31:0] local_bb2_shl273_i604;

assign local_bb2_shl273_i604 = (rnode_189to190_bb2_and269_i603_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp258_i597_stall_local;
wire local_bb2_cmp258_i597;

assign local_bb2_cmp258_i597 = ($signed(rnode_189to190_bb2_add245_i589_0_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb2_and272_i602_stall_local;
wire [31:0] local_bb2_and272_i602;

assign local_bb2_and272_i602 = (rnode_189to190_bb2_shr271_i601_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp226_not_i584_stall_local;
wire local_bb2_cmp226_not_i584;

assign local_bb2_cmp226_not_i584 = (rnode_189to190_bb2_cmp226_i583_0_NO_SHIFT_REG ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb2__47_i596_stall_local;
wire local_bb2__47_i596;

assign local_bb2__47_i596 = (rnode_189to190_bb2_cmp226_i583_1_NO_SHIFT_REG | rnode_189to190_bb2_not__46_i595_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp29649_i619_stall_local;
wire [31:0] local_bb2_cmp29649_i619;

assign local_bb2_cmp29649_i619[31:1] = 31'h0;
assign local_bb2_cmp29649_i619[0] = rnode_189to190_bb2_cmp296_i615_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_conv300_i617_stall_local;
wire [31:0] local_bb2_conv300_i617;

assign local_bb2_conv300_i617[31:1] = 31'h0;
assign local_bb2_conv300_i617[0] = rnode_189to190_bb2_cmp299_i616_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_shl273_i_stall_local;
wire [31:0] local_bb2_shl273_i;

assign local_bb2_shl273_i = (rnode_189to190_bb2_and269_i_0_NO_SHIFT_REG & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb2_cmp258_i_stall_local;
wire local_bb2_cmp258_i;

assign local_bb2_cmp258_i = ($signed(rnode_189to190_bb2_add245_i_0_NO_SHIFT_REG) > $signed(32'hFE));

// This section implements an unregistered operation.
// 
wire local_bb2_and272_i_stall_local;
wire [31:0] local_bb2_and272_i;

assign local_bb2_and272_i = (rnode_189to190_bb2_shr271_i_0_NO_SHIFT_REG & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u170_valid_out;
wire local_bb2_var__u170_stall_in;
wire local_bb2_var__u170_inputs_ready;
wire local_bb2_var__u170_stall_local;
wire [31:0] local_bb2_var__u170;

assign local_bb2_var__u170_inputs_ready = rnode_189to190_bb2__47_i_0_valid_out_1_NO_SHIFT_REG;
assign local_bb2_var__u170[31:1] = 31'h0;
assign local_bb2_var__u170[0] = rnode_189to190_bb2__47_i_1_NO_SHIFT_REG;
assign local_bb2_var__u170_valid_out = 1'b1;
assign rnode_189to190_bb2__47_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;

// This section implements an unregistered operation.
// 
wire local_bb2_cmp29649_i_stall_local;
wire [31:0] local_bb2_cmp29649_i;

assign local_bb2_cmp29649_i[31:1] = 31'h0;
assign local_bb2_cmp29649_i[0] = rnode_189to190_bb2_cmp296_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_conv300_i_stall_local;
wire [31:0] local_bb2_conv300_i;

assign local_bb2_conv300_i[31:1] = 31'h0;
assign local_bb2_conv300_i[0] = rnode_189to190_bb2_cmp299_i_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge12_i_stall_local;
wire local_bb2_brmerge12_i;

assign local_bb2_brmerge12_i = (rnode_189to190_bb2_cmp226_not_i_0_NO_SHIFT_REG | rnode_189to190_bb2_not_cmp37_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_or274_i605_stall_local;
wire [31:0] local_bb2_or274_i605;

assign local_bb2_or274_i605 = (local_bb2_and272_i602 | local_bb2_shl273_i604);

// This section implements an unregistered operation.
// 
wire local_bb2_brmerge12_i585_stall_local;
wire local_bb2_brmerge12_i585;

assign local_bb2_brmerge12_i585 = (local_bb2_cmp226_not_i584 | rnode_189to190_bb2_not_cmp37_i577_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot262__i598_stall_local;
wire local_bb2_lnot262__i598;

assign local_bb2_lnot262__i598 = (local_bb2_cmp258_i597 & local_bb2_cmp226_not_i584);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot262__i_stall_local;
wire local_bb2_lnot262__i;

assign local_bb2_lnot262__i = (local_bb2_cmp258_i & rnode_189to190_bb2_cmp226_not_i_1_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_or274_i_stall_local;
wire [31:0] local_bb2_or274_i;

assign local_bb2_or274_i = (local_bb2_and272_i | local_bb2_shl273_i);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_var__u170_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_var__u170_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_var__u170_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_var__u170_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_var__u170_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_var__u170_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_var__u170_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_var__u170_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_var__u170_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_var__u170_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_var__u170_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_var__u170_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_var__u170_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(local_bb2_var__u170),
	.data_out(rnode_190to191_bb2_var__u170_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_var__u170_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_var__u170_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_var__u170_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_var__u170_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_var__u170_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_var__u170_stall_in = 1'b0;
assign rnode_190to191_bb2_var__u170_0_NO_SHIFT_REG = rnode_190to191_bb2_var__u170_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_var__u170_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_var__u170_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_resultSign_0_i_stall_local;
wire [31:0] local_bb2_resultSign_0_i;

assign local_bb2_resultSign_0_i = (local_bb2_brmerge12_i ? rnode_189to190_bb2_and35_i_0_NO_SHIFT_REG : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_resultSign_0_i586_stall_local;
wire [31:0] local_bb2_resultSign_0_i586;

assign local_bb2_resultSign_0_i586 = (local_bb2_brmerge12_i585 ? rnode_189to190_bb2_and35_i469_0_NO_SHIFT_REG : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_or2662_i599_stall_local;
wire local_bb2_or2662_i599;

assign local_bb2_or2662_i599 = (rnode_189to190_bb2_var__u157_0_NO_SHIFT_REG | local_bb2_lnot262__i598);

// This section implements an unregistered operation.
// 
wire local_bb2_or2662_i_stall_local;
wire local_bb2_or2662_i;

assign local_bb2_or2662_i = (rnode_189to190_bb2_var__u156_0_NO_SHIFT_REG | local_bb2_lnot262__i);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext314_i_stall_local;
wire [31:0] local_bb2_lnot_ext314_i;

assign local_bb2_lnot_ext314_i = (rnode_190to191_bb2_var__u170_0_NO_SHIFT_REG ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_or275_i_stall_local;
wire [31:0] local_bb2_or275_i;

assign local_bb2_or275_i = (local_bb2_or274_i | local_bb2_resultSign_0_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or275_i606_stall_local;
wire [31:0] local_bb2_or275_i606;

assign local_bb2_or275_i606 = (local_bb2_or274_i605 | local_bb2_resultSign_0_i586);

// This section implements an unregistered operation.
// 
wire local_bb2_or2804_i607_stall_local;
wire local_bb2_or2804_i607;

assign local_bb2_or2804_i607 = (local_bb2__47_i596 | local_bb2_or2662_i599);

// This section implements an unregistered operation.
// 
wire local_bb2_or2875_i609_stall_local;
wire local_bb2_or2875_i609;

assign local_bb2_or2875_i609 = (local_bb2_or2662_i599 | rnode_189to190_bb2__26_i484_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u171_stall_local;
wire [31:0] local_bb2_var__u171;

assign local_bb2_var__u171[31:1] = 31'h0;
assign local_bb2_var__u171[0] = local_bb2_or2662_i599;

// This section implements an unregistered operation.
// 
wire local_bb2_or2804_i_stall_local;
wire local_bb2_or2804_i;

assign local_bb2_or2804_i = (rnode_189to190_bb2__47_i_0_NO_SHIFT_REG | local_bb2_or2662_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or2875_i_stall_local;
wire local_bb2_or2875_i;

assign local_bb2_or2875_i = (local_bb2_or2662_i | rnode_189to190_bb2__26_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u172_stall_local;
wire [31:0] local_bb2_var__u172;

assign local_bb2_var__u172[31:1] = 31'h0;
assign local_bb2_var__u172[0] = local_bb2_or2662_i;

// This section implements an unregistered operation.
// 
wire local_bb2_cond282_i608_stall_local;
wire [31:0] local_bb2_cond282_i608;

assign local_bb2_cond282_i608 = (local_bb2_or2804_i607 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond289_i610_stall_local;
wire [31:0] local_bb2_cond289_i610;

assign local_bb2_cond289_i610 = (local_bb2_or2875_i609 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext310_i622_stall_local;
wire [31:0] local_bb2_lnot_ext310_i622;

assign local_bb2_lnot_ext310_i622 = (local_bb2_var__u171 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_cond282_i_stall_local;
wire [31:0] local_bb2_cond282_i;

assign local_bb2_cond282_i = (local_bb2_or2804_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb2_cond289_i_stall_local;
wire [31:0] local_bb2_cond289_i;

assign local_bb2_cond289_i = (local_bb2_or2875_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext310_i_stall_local;
wire [31:0] local_bb2_lnot_ext310_i;

assign local_bb2_lnot_ext310_i = (local_bb2_var__u172 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_and293_i612_stall_local;
wire [31:0] local_bb2_and293_i612;

assign local_bb2_and293_i612 = (local_bb2_cond282_i608 & local_bb2_or275_i606);

// This section implements an unregistered operation.
// 
wire local_bb2_or294_i613_stall_local;
wire [31:0] local_bb2_or294_i613;

assign local_bb2_or294_i613 = (local_bb2_cond289_i610 | local_bb2_cond292_i611);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i624_stall_local;
wire [31:0] local_bb2_reduction_0_i624;

assign local_bb2_reduction_0_i624 = (local_bb2_lnot_ext310_i622 & local_bb2_lnot_ext_i621);

// This section implements an unregistered operation.
// 
wire local_bb2_and293_i_stall_local;
wire [31:0] local_bb2_and293_i;

assign local_bb2_and293_i = (local_bb2_cond282_i & local_bb2_or275_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or294_i_stall_local;
wire [31:0] local_bb2_or294_i;

assign local_bb2_or294_i = (local_bb2_cond289_i | local_bb2_cond292_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_0_i78_stall_local;
wire [31:0] local_bb2_reduction_0_i78;

assign local_bb2_reduction_0_i78 = (local_bb2_lnot_ext310_i & local_bb2_lnot_ext_i);

// This section implements an unregistered operation.
// 
wire local_bb2_and302_i618_stall_local;
wire [31:0] local_bb2_and302_i618;

assign local_bb2_and302_i618 = (local_bb2_conv300_i617 & local_bb2_and293_i612);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i614_stall_local;
wire [31:0] local_bb2_or295_i614;

assign local_bb2_or295_i614 = (local_bb2_or294_i613 | local_bb2_and293_i612);

// This section implements an unregistered operation.
// 
wire local_bb2_and302_i_stall_local;
wire [31:0] local_bb2_and302_i;

assign local_bb2_and302_i = (local_bb2_conv300_i & local_bb2_and293_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i_stall_local;
wire [31:0] local_bb2_or295_i;

assign local_bb2_or295_i = (local_bb2_or294_i | local_bb2_and293_i);

// This section implements an unregistered operation.
// 
wire local_bb2_or295_i614_valid_out;
wire local_bb2_or295_i614_stall_in;
 reg local_bb2_or295_i614_consumed_0_NO_SHIFT_REG;
wire local_bb2__47_i596_valid_out_1;
wire local_bb2__47_i596_stall_in_1;
 reg local_bb2__47_i596_consumed_1_NO_SHIFT_REG;
wire local_bb2_lor_ext_i620_valid_out;
wire local_bb2_lor_ext_i620_stall_in;
 reg local_bb2_lor_ext_i620_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i624_valid_out;
wire local_bb2_reduction_0_i624_stall_in;
 reg local_bb2_reduction_0_i624_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i620_inputs_ready;
wire local_bb2_lor_ext_i620_stall_local;
wire [31:0] local_bb2_lor_ext_i620;

assign local_bb2_lor_ext_i620_inputs_ready = (rnode_189to190_bb2_and35_i469_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_not_cmp37_i577_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_and269_i603_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_add245_i589_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_var__u157_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2__26_i484_0_valid_out_0_NO_SHIFT_REG & rnode_189to190_bb2__26_i484_0_valid_out_1_NO_SHIFT_REG & rnode_189to190_bb2_cmp226_i583_0_valid_out_1_NO_SHIFT_REG & rnode_189to190_bb2_not__46_i595_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_shr271_i601_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2__26_i484_0_valid_out_2_NO_SHIFT_REG & rnode_189to190_bb2_cmp226_i583_0_valid_out_0_NO_SHIFT_REG & rnode_189to190_bb2_cmp296_i615_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_cmp299_i616_0_valid_out_NO_SHIFT_REG);
assign local_bb2_lor_ext_i620 = (local_bb2_cmp29649_i619 | local_bb2_and302_i618);
assign local_bb2_or295_i614_valid_out = 1'b1;
assign local_bb2__47_i596_valid_out_1 = 1'b1;
assign local_bb2_lor_ext_i620_valid_out = 1'b1;
assign local_bb2_reduction_0_i624_valid_out = 1'b1;
assign rnode_189to190_bb2_and35_i469_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_not_cmp37_i577_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_and269_i603_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_add245_i589_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_var__u157_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i484_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i484_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp226_i583_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_not__46_i595_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_shr271_i601_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i484_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp226_i583_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp296_i615_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp299_i616_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_or295_i614_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2__47_i596_consumed_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_lor_ext_i620_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i624_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_or295_i614_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i620_inputs_ready & (local_bb2_or295_i614_consumed_0_NO_SHIFT_REG | ~(local_bb2_or295_i614_stall_in)) & local_bb2_lor_ext_i620_stall_local);
		local_bb2__47_i596_consumed_1_NO_SHIFT_REG <= (local_bb2_lor_ext_i620_inputs_ready & (local_bb2__47_i596_consumed_1_NO_SHIFT_REG | ~(local_bb2__47_i596_stall_in_1)) & local_bb2_lor_ext_i620_stall_local);
		local_bb2_lor_ext_i620_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i620_inputs_ready & (local_bb2_lor_ext_i620_consumed_0_NO_SHIFT_REG | ~(local_bb2_lor_ext_i620_stall_in)) & local_bb2_lor_ext_i620_stall_local);
		local_bb2_reduction_0_i624_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i620_inputs_ready & (local_bb2_reduction_0_i624_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i624_stall_in)) & local_bb2_lor_ext_i620_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_or295_i_valid_out;
wire local_bb2_or295_i_stall_in;
 reg local_bb2_or295_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i_valid_out;
wire local_bb2_lor_ext_i_stall_in;
 reg local_bb2_lor_ext_i_consumed_0_NO_SHIFT_REG;
wire local_bb2_reduction_0_i78_valid_out;
wire local_bb2_reduction_0_i78_stall_in;
 reg local_bb2_reduction_0_i78_consumed_0_NO_SHIFT_REG;
wire local_bb2_lor_ext_i_inputs_ready;
wire local_bb2_lor_ext_i_stall_local;
wire [31:0] local_bb2_lor_ext_i;

assign local_bb2_lor_ext_i_inputs_ready = (rnode_189to190_bb2_and35_i_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_cmp226_not_i_0_valid_out_0_NO_SHIFT_REG & rnode_189to190_bb2_not_cmp37_i_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_and269_i_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_add245_i_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_cmp226_not_i_0_valid_out_1_NO_SHIFT_REG & rnode_189to190_bb2_var__u156_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2__47_i_0_valid_out_0_NO_SHIFT_REG & rnode_189to190_bb2__26_i_0_valid_out_0_NO_SHIFT_REG & rnode_189to190_bb2__26_i_0_valid_out_1_NO_SHIFT_REG & rnode_189to190_bb2_shr271_i_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2__26_i_0_valid_out_2_NO_SHIFT_REG & rnode_189to190_bb2_cmp296_i_0_valid_out_NO_SHIFT_REG & rnode_189to190_bb2_cmp299_i_0_valid_out_NO_SHIFT_REG);
assign local_bb2_lor_ext_i = (local_bb2_cmp29649_i | local_bb2_and302_i);
assign local_bb2_or295_i_valid_out = 1'b1;
assign local_bb2_lor_ext_i_valid_out = 1'b1;
assign local_bb2_reduction_0_i78_valid_out = 1'b1;
assign rnode_189to190_bb2_and35_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp226_not_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_not_cmp37_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_and269_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_add245_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp226_not_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_var__u156_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__47_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i_0_stall_in_0_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i_0_stall_in_1_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_shr271_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2__26_i_0_stall_in_2_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp296_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_189to190_bb2_cmp299_i_0_stall_in_NO_SHIFT_REG = 1'b0;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_or295_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_lor_ext_i_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_reduction_0_i78_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_or295_i_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i_inputs_ready & (local_bb2_or295_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_or295_i_stall_in)) & local_bb2_lor_ext_i_stall_local);
		local_bb2_lor_ext_i_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i_inputs_ready & (local_bb2_lor_ext_i_consumed_0_NO_SHIFT_REG | ~(local_bb2_lor_ext_i_stall_in)) & local_bb2_lor_ext_i_stall_local);
		local_bb2_reduction_0_i78_consumed_0_NO_SHIFT_REG <= (local_bb2_lor_ext_i_inputs_ready & (local_bb2_reduction_0_i78_consumed_0_NO_SHIFT_REG | ~(local_bb2_reduction_0_i78_stall_in)) & local_bb2_lor_ext_i_stall_local);
	end
end


// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_or295_i614_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i614_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_or295_i614_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i614_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_or295_i614_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i614_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i614_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i614_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_or295_i614_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_or295_i614_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_or295_i614_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_or295_i614_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_or295_i614_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(local_bb2_or295_i614),
	.data_out(rnode_190to191_bb2_or295_i614_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_or295_i614_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_or295_i614_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_or295_i614_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_or295_i614_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_or295_i614_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or295_i614_stall_in = 1'b0;
assign rnode_190to191_bb2_or295_i614_0_NO_SHIFT_REG = rnode_190to191_bb2_or295_i614_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_or295_i614_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_or295_i614_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2__47_i596_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2__47_i596_0_stall_in_NO_SHIFT_REG;
 logic rnode_190to191_bb2__47_i596_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2__47_i596_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic rnode_190to191_bb2__47_i596_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2__47_i596_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2__47_i596_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2__47_i596_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2__47_i596_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2__47_i596_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2__47_i596_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2__47_i596_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2__47_i596_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(local_bb2__47_i596),
	.data_out(rnode_190to191_bb2__47_i596_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2__47_i596_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2__47_i596_0_reg_191_fifo.DATA_WIDTH = 1;
defparam rnode_190to191_bb2__47_i596_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2__47_i596_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2__47_i596_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2__47_i596_stall_in_1 = 1'b0;
assign rnode_190to191_bb2__47_i596_0_NO_SHIFT_REG = rnode_190to191_bb2__47_i596_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2__47_i596_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2__47_i596_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_lor_ext_i620_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i620_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_lor_ext_i620_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i620_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_lor_ext_i620_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i620_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i620_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i620_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_lor_ext_i620_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_lor_ext_i620_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_lor_ext_i620_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_lor_ext_i620_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_lor_ext_i620_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(local_bb2_lor_ext_i620),
	.data_out(rnode_190to191_bb2_lor_ext_i620_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_lor_ext_i620_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_lor_ext_i620_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_lor_ext_i620_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_lor_ext_i620_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_lor_ext_i620_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lor_ext_i620_stall_in = 1'b0;
assign rnode_190to191_bb2_lor_ext_i620_0_NO_SHIFT_REG = rnode_190to191_bb2_lor_ext_i620_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_lor_ext_i620_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_lor_ext_i620_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_reduction_0_i624_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i624_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_reduction_0_i624_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i624_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_reduction_0_i624_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i624_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i624_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i624_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_reduction_0_i624_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_reduction_0_i624_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_reduction_0_i624_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_reduction_0_i624_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_reduction_0_i624_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i624),
	.data_out(rnode_190to191_bb2_reduction_0_i624_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_reduction_0_i624_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_reduction_0_i624_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_reduction_0_i624_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_reduction_0_i624_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_reduction_0_i624_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i624_stall_in = 1'b0;
assign rnode_190to191_bb2_reduction_0_i624_0_NO_SHIFT_REG = rnode_190to191_bb2_reduction_0_i624_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_reduction_0_i624_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_reduction_0_i624_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_or295_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_or295_i_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_or295_i_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_or295_i_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_or295_i_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_or295_i_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_or295_i_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_or295_i_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_or295_i_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(local_bb2_or295_i),
	.data_out(rnode_190to191_bb2_or295_i_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_or295_i_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_or295_i_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_or295_i_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_or295_i_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_or295_i_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_or295_i_stall_in = 1'b0;
assign rnode_190to191_bb2_or295_i_0_NO_SHIFT_REG = rnode_190to191_bb2_or295_i_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_or295_i_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_or295_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_lor_ext_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_lor_ext_i_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_lor_ext_i_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_lor_ext_i_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_lor_ext_i_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_lor_ext_i_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_lor_ext_i_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_lor_ext_i_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_lor_ext_i_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(local_bb2_lor_ext_i),
	.data_out(rnode_190to191_bb2_lor_ext_i_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_lor_ext_i_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_lor_ext_i_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_lor_ext_i_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_lor_ext_i_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_lor_ext_i_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_lor_ext_i_stall_in = 1'b0;
assign rnode_190to191_bb2_lor_ext_i_0_NO_SHIFT_REG = rnode_190to191_bb2_lor_ext_i_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_lor_ext_i_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_lor_ext_i_0_valid_out_NO_SHIFT_REG = 1'b1;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_190to191_bb2_reduction_0_i78_0_valid_out_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i78_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_reduction_0_i78_0_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i78_0_reg_191_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_190to191_bb2_reduction_0_i78_0_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i78_0_valid_out_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i78_0_stall_in_reg_191_NO_SHIFT_REG;
 logic rnode_190to191_bb2_reduction_0_i78_0_stall_out_reg_191_NO_SHIFT_REG;

acl_data_fifo rnode_190to191_bb2_reduction_0_i78_0_reg_191_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_190to191_bb2_reduction_0_i78_0_reg_191_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_190to191_bb2_reduction_0_i78_0_stall_in_reg_191_NO_SHIFT_REG),
	.valid_out(rnode_190to191_bb2_reduction_0_i78_0_valid_out_reg_191_NO_SHIFT_REG),
	.stall_out(rnode_190to191_bb2_reduction_0_i78_0_stall_out_reg_191_NO_SHIFT_REG),
	.data_in(local_bb2_reduction_0_i78),
	.data_out(rnode_190to191_bb2_reduction_0_i78_0_reg_191_NO_SHIFT_REG)
);

defparam rnode_190to191_bb2_reduction_0_i78_0_reg_191_fifo.DEPTH = 1;
defparam rnode_190to191_bb2_reduction_0_i78_0_reg_191_fifo.DATA_WIDTH = 32;
defparam rnode_190to191_bb2_reduction_0_i78_0_reg_191_fifo.ALLOW_FULL_WRITE = 1;
defparam rnode_190to191_bb2_reduction_0_i78_0_reg_191_fifo.IMPL = "shift_reg";

assign rnode_190to191_bb2_reduction_0_i78_0_reg_191_inputs_ready_NO_SHIFT_REG = 1'b1;
assign local_bb2_reduction_0_i78_stall_in = 1'b0;
assign rnode_190to191_bb2_reduction_0_i78_0_NO_SHIFT_REG = rnode_190to191_bb2_reduction_0_i78_0_reg_191_NO_SHIFT_REG;
assign rnode_190to191_bb2_reduction_0_i78_0_stall_in_reg_191_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_reduction_0_i78_0_valid_out_NO_SHIFT_REG = 1'b1;

// This section implements an unregistered operation.
// 
wire local_bb2_var__u173_stall_local;
wire [31:0] local_bb2_var__u173;

assign local_bb2_var__u173[31:1] = 31'h0;
assign local_bb2_var__u173[0] = rnode_190to191_bb2__47_i596_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_1_i_stall_local;
wire [31:0] local_bb2_reduction_1_i;

assign local_bb2_reduction_1_i = (local_bb2_lnot_ext314_i & rnode_190to191_bb2_lor_ext_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_lnot_ext314_i623_stall_local;
wire [31:0] local_bb2_lnot_ext314_i623;

assign local_bb2_lnot_ext314_i623 = (local_bb2_var__u173 ^ 32'h1);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i79_stall_local;
wire [31:0] local_bb2_reduction_2_i79;

assign local_bb2_reduction_2_i79 = (rnode_190to191_bb2_reduction_0_i78_0_NO_SHIFT_REG & local_bb2_reduction_1_i);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_1_i625_stall_local;
wire [31:0] local_bb2_reduction_1_i625;

assign local_bb2_reduction_1_i625 = (local_bb2_lnot_ext314_i623 & rnode_190to191_bb2_lor_ext_i620_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_add320_i_stall_local;
wire [31:0] local_bb2_add320_i;

assign local_bb2_add320_i = (local_bb2_reduction_2_i79 + rnode_190to191_bb2_or295_i_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_reduction_2_i626_stall_local;
wire [31:0] local_bb2_reduction_2_i626;

assign local_bb2_reduction_2_i626 = (rnode_190to191_bb2_reduction_0_i624_0_NO_SHIFT_REG & local_bb2_reduction_1_i625);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u174_stall_local;
wire [31:0] local_bb2_var__u174;

assign local_bb2_var__u174 = local_bb2_add320_i;

// This section implements an unregistered operation.
// 
wire local_bb2_add320_i627_stall_local;
wire [31:0] local_bb2_add320_i627;

assign local_bb2_add320_i627 = (local_bb2_reduction_2_i626 + rnode_190to191_bb2_or295_i614_0_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb2_var__u175_stall_local;
wire [31:0] local_bb2_var__u175;

assign local_bb2_var__u175 = local_bb2_add320_i627;

// This section implements an unregistered operation.
// 
wire local_bb2_c0_exi3_stall_local;
wire [159:0] local_bb2_c0_exi3;

assign local_bb2_c0_exi3[95:0] = local_bb2_c0_exi2[95:0];
assign local_bb2_c0_exi3[127:96] = local_bb2_var__u175;
assign local_bb2_c0_exi3[159:128] = local_bb2_c0_exi2[159:128];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_exi4_valid_out;
wire local_bb2_c0_exi4_stall_in;
wire local_bb2_c0_exi4_inputs_ready;
wire local_bb2_c0_exi4_stall_local;
wire [159:0] local_bb2_c0_exi4;

assign local_bb2_c0_exi4_inputs_ready = (rnode_190to191_bb2_add320_i1639_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2_add320_i1091_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2_or295_i614_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2_reduction_0_i624_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2__47_i596_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2_lor_ext_i620_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2_or295_i_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2_reduction_0_i78_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2_var__u170_0_valid_out_NO_SHIFT_REG & rnode_190to191_bb2_lor_ext_i_0_valid_out_NO_SHIFT_REG);
assign local_bb2_c0_exi4[127:0] = local_bb2_c0_exi3[127:0];
assign local_bb2_c0_exi4[159:128] = local_bb2_var__u174;
assign local_bb2_c0_exi4_valid_out = 1'b1;
assign rnode_190to191_bb2_add320_i1639_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_add320_i1091_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_or295_i614_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_reduction_0_i624_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2__47_i596_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_lor_ext_i620_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_or295_i_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_reduction_0_i78_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_var__u170_0_stall_in_NO_SHIFT_REG = 1'b0;
assign rnode_190to191_bb2_lor_ext_i_0_stall_in_NO_SHIFT_REG = 1'b0;

// This section implements a registered operation.
// 
wire local_bb2_c0_exit_c0_exi4_inputs_ready;
 reg local_bb2_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG;
wire local_bb2_c0_exit_c0_exi4_stall_in_0;
 reg local_bb2_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG;
wire local_bb2_c0_exit_c0_exi4_stall_in_1;
 reg local_bb2_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG;
wire local_bb2_c0_exit_c0_exi4_stall_in_2;
 reg [159:0] local_bb2_c0_exit_c0_exi4_NO_SHIFT_REG;
wire [159:0] local_bb2_c0_exit_c0_exi4_in;
wire local_bb2_c0_exit_c0_exi4_valid;
wire local_bb2_c0_exit_c0_exi4_causedstall;

acl_stall_free_sink local_bb2_c0_exit_c0_exi4_instance (
	.clock(clock),
	.resetn(resetn),
	.data_in(local_bb2_c0_exi4),
	.data_out(local_bb2_c0_exit_c0_exi4_in),
	.input_accepted(local_bb2_c0_enter_c0_eni8_input_accepted),
	.valid_out(local_bb2_c0_exit_c0_exi4_valid),
	.stall_in(~(local_bb2_c0_exit_c0_exi4_output_regs_ready)),
	.stall_entry(local_bb2_c0_exit_c0_exi4_entry_stall),
	.valids(local_bb2_c0_exit_c0_exi4_valid_bits),
	.IIphases(local_bb2_c0_exit_c0_exi4_phases),
	.inc_pipelined_thread(local_bb2_c0_enter_c0_eni8_inc_pipelined_thread),
	.dec_pipelined_thread(local_bb2_c0_enter_c0_eni8_dec_pipelined_thread)
);

defparam local_bb2_c0_exit_c0_exi4_instance.DATA_WIDTH = 160;
defparam local_bb2_c0_exit_c0_exi4_instance.PIPELINE_DEPTH = 31;
defparam local_bb2_c0_exit_c0_exi4_instance.SHARINGII = 1;
defparam local_bb2_c0_exit_c0_exi4_instance.SCHEDULEII = 1;

assign local_bb2_c0_exit_c0_exi4_inputs_ready = 1'b1;
assign local_bb2_c0_exit_c0_exi4_output_regs_ready = ((~(local_bb2_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG) | ~(local_bb2_c0_exit_c0_exi4_stall_in_0)) & (~(local_bb2_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG) | ~(local_bb2_c0_exit_c0_exi4_stall_in_1)) & (~(local_bb2_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG) | ~(local_bb2_c0_exit_c0_exi4_stall_in_2)));
assign local_bb2_c0_exi4_stall_in = 1'b0;
assign local_bb2_c0_exit_c0_exi4_causedstall = (1'b1 && (1'b0 && !(~(local_bb2_c0_exit_c0_exi4_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_c0_exit_c0_exi4_NO_SHIFT_REG <= 'x;
		local_bb2_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb2_c0_exit_c0_exi4_output_regs_ready)
		begin
			local_bb2_c0_exit_c0_exi4_NO_SHIFT_REG <= local_bb2_c0_exit_c0_exi4_in;
			local_bb2_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= local_bb2_c0_exit_c0_exi4_valid;
			local_bb2_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= local_bb2_c0_exit_c0_exi4_valid;
			local_bb2_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= local_bb2_c0_exit_c0_exi4_valid;
		end
		else
		begin
			if (~(local_bb2_c0_exit_c0_exi4_stall_in_0))
			begin
				local_bb2_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_exit_c0_exi4_stall_in_1))
			begin
				local_bb2_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(local_bb2_c0_exit_c0_exi4_stall_in_2))
			begin
				local_bb2_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements an unregistered operation.
// 
wire local_bb2_c0_exe3_stall_local;
wire [31:0] local_bb2_c0_exe3;

assign local_bb2_c0_exe3 = local_bb2_c0_exit_c0_exi4_NO_SHIFT_REG[127:96];

// This section implements an unregistered operation.
// 
wire local_bb2_c0_exe4_valid_out;
wire local_bb2_c0_exe4_stall_in;
 reg local_bb2_c0_exe4_consumed_0_NO_SHIFT_REG;
wire local_bb2_c0_exe3_valid_out;
wire local_bb2_c0_exe3_stall_in;
 reg local_bb2_c0_exe3_consumed_0_NO_SHIFT_REG;
wire local_bb2_c0_exe4_inputs_ready;
wire local_bb2_c0_exe4_stall_local;
wire [31:0] local_bb2_c0_exe4;

assign local_bb2_c0_exe4_inputs_ready = (local_bb2_c0_exit_c0_exi4_valid_out_1_NO_SHIFT_REG & local_bb2_c0_exit_c0_exi4_valid_out_0_NO_SHIFT_REG);
assign local_bb2_c0_exe4 = local_bb2_c0_exit_c0_exi4_NO_SHIFT_REG[159:128];
assign local_bb2_c0_exe4_stall_local = ((local_bb2_c0_exe4_stall_in & ~(local_bb2_c0_exe4_consumed_0_NO_SHIFT_REG)) | (local_bb2_c0_exe3_stall_in & ~(local_bb2_c0_exe3_consumed_0_NO_SHIFT_REG)));
assign local_bb2_c0_exe4_valid_out = (local_bb2_c0_exe4_inputs_ready & ~(local_bb2_c0_exe4_consumed_0_NO_SHIFT_REG));
assign local_bb2_c0_exe3_valid_out = (local_bb2_c0_exe4_inputs_ready & ~(local_bb2_c0_exe3_consumed_0_NO_SHIFT_REG));
assign local_bb2_c0_exit_c0_exi4_stall_in_1 = (local_bb2_c0_exe4_stall_local | ~(local_bb2_c0_exe4_inputs_ready));
assign local_bb2_c0_exit_c0_exi4_stall_in_0 = (local_bb2_c0_exe4_stall_local | ~(local_bb2_c0_exe4_inputs_ready));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb2_c0_exe4_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb2_c0_exe3_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb2_c0_exe4_consumed_0_NO_SHIFT_REG <= (local_bb2_c0_exe4_inputs_ready & (local_bb2_c0_exe4_consumed_0_NO_SHIFT_REG | ~(local_bb2_c0_exe4_stall_in)) & local_bb2_c0_exe4_stall_local);
		local_bb2_c0_exe3_consumed_0_NO_SHIFT_REG <= (local_bb2_c0_exe4_inputs_ready & (local_bb2_c0_exe3_consumed_0_NO_SHIFT_REG | ~(local_bb2_c0_exe3_stall_in)) & local_bb2_c0_exe4_stall_local);
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
 reg branch_node_valid_out_0_NO_SHIFT_REG;
 reg branch_compare_result_NO_SHIFT_REG;
wire branch_var__output_regs_ready;
wire combined_branch_stall_in_signal;
 reg [63:0] lvb_var__0_reg_NO_SHIFT_REG;
 reg [63:0] lvb_bb2_indvars_iv_next_1_0_reg_NO_SHIFT_REG;
 reg lvb_bb2_exitcond_0_reg_NO_SHIFT_REG;
 reg [159:0] lvb_bb2_c0_exit_c0_exi4_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb2_c0_exe3_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_bb2_c0_exe4_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
 reg [31:0] lvb_input_global_id_1_0_reg_NO_SHIFT_REG;

assign branch_var__inputs_ready = (local_bb2_c0_exe4_valid_out & local_bb2_c0_exe3_valid_out & local_bb2__24_demorgan_GUARD_valid_out & local_bb2_c0_exit_c0_exi4_valid_out_2_NO_SHIFT_REG & rnode_195to196_bb2_indvars_iv_next_1_0_valid_out_1_NO_SHIFT_REG & rnode_195to196_input_global_id_1_0_valid_out_NO_SHIFT_REG & rnode_195to196_var__0_valid_out_NO_SHIFT_REG & rnode_195to196_input_global_id_0_0_valid_out_NO_SHIFT_REG & rnode_195to196_bb2_exitcond_0_valid_out_1_NO_SHIFT_REG);
assign branch_var__output_regs_ready = (~(branch_node_valid_out_0_NO_SHIFT_REG) | (((branch_compare_result_NO_SHIFT_REG != 1'b1) & ~(stall_in_1)) | (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & ~(stall_in_0))));
assign local_bb2_c0_exe4_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb2_c0_exe3_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb2__24_demorgan_GUARD_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign local_bb2_c0_exit_c0_exi4_stall_in_2 = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_195to196_bb2_indvars_iv_next_1_0_stall_in_1_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_195to196_input_global_id_1_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_195to196_var__0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_195to196_input_global_id_0_0_stall_in_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign rnode_195to196_bb2_exitcond_0_stall_in_1_NO_SHIFT_REG = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign lvb_var__0 = lvb_var__0_reg_NO_SHIFT_REG;
assign lvb_var__1 = lvb_var__0_reg_NO_SHIFT_REG;
assign lvb_bb2_indvars_iv_next_1_0 = lvb_bb2_indvars_iv_next_1_0_reg_NO_SHIFT_REG;
assign lvb_bb2_indvars_iv_next_1_1 = lvb_bb2_indvars_iv_next_1_0_reg_NO_SHIFT_REG;
assign lvb_bb2_exitcond_0 = lvb_bb2_exitcond_0_reg_NO_SHIFT_REG;
assign lvb_bb2_exitcond_1 = lvb_bb2_exitcond_0_reg_NO_SHIFT_REG;
assign lvb_bb2_c0_exit_c0_exi4_0 = lvb_bb2_c0_exit_c0_exi4_0_reg_NO_SHIFT_REG;
assign lvb_bb2_c0_exit_c0_exi4_1 = lvb_bb2_c0_exit_c0_exi4_0_reg_NO_SHIFT_REG;
assign lvb_bb2_c0_exe3_0 = lvb_bb2_c0_exe3_0_reg_NO_SHIFT_REG;
assign lvb_bb2_c0_exe3_1 = lvb_bb2_c0_exe3_0_reg_NO_SHIFT_REG;
assign lvb_bb2_c0_exe4_0 = lvb_bb2_c0_exe4_0_reg_NO_SHIFT_REG;
assign lvb_bb2_c0_exe4_1 = lvb_bb2_c0_exe4_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0_0 = lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_0_1 = lvb_input_global_id_0_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1_0 = lvb_input_global_id_1_0_reg_NO_SHIFT_REG;
assign lvb_input_global_id_1_1 = lvb_input_global_id_1_0_reg_NO_SHIFT_REG;
assign valid_out_0 = (~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG);
assign valid_out_1 = ((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG);
assign combined_branch_stall_in_signal = ((((branch_compare_result_NO_SHIFT_REG != 1'b1) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_1) | ((~((branch_compare_result_NO_SHIFT_REG != 1'b1)) & branch_node_valid_out_0_NO_SHIFT_REG) & stall_in_0));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		lvb_var__0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_indvars_iv_next_1_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_exitcond_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_c0_exit_c0_exi4_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_c0_exe3_0_reg_NO_SHIFT_REG <= 'x;
		lvb_bb2_c0_exe4_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_0_0_reg_NO_SHIFT_REG <= 'x;
		lvb_input_global_id_1_0_reg_NO_SHIFT_REG <= 'x;
		branch_compare_result_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (branch_var__output_regs_ready)
		begin
			branch_node_valid_out_0_NO_SHIFT_REG <= branch_var__inputs_ready;
			lvb_var__0_reg_NO_SHIFT_REG <= rnode_195to196_var__0_NO_SHIFT_REG;
			lvb_bb2_indvars_iv_next_1_0_reg_NO_SHIFT_REG <= rnode_195to196_bb2_indvars_iv_next_1_1_NO_SHIFT_REG;
			lvb_bb2_exitcond_0_reg_NO_SHIFT_REG <= rnode_195to196_bb2_exitcond_1_NO_SHIFT_REG;
			lvb_bb2_c0_exit_c0_exi4_0_reg_NO_SHIFT_REG <= local_bb2_c0_exit_c0_exi4_NO_SHIFT_REG;
			lvb_bb2_c0_exe3_0_reg_NO_SHIFT_REG <= local_bb2_c0_exe3;
			lvb_bb2_c0_exe4_0_reg_NO_SHIFT_REG <= local_bb2_c0_exe4;
			lvb_input_global_id_0_0_reg_NO_SHIFT_REG <= rnode_195to196_input_global_id_0_0_NO_SHIFT_REG;
			lvb_input_global_id_1_0_reg_NO_SHIFT_REG <= rnode_195to196_input_global_id_1_0_NO_SHIFT_REG;
			branch_compare_result_NO_SHIFT_REG <= local_bb2__24_demorgan_GUARD;
		end
		else
		begin
			if (~(combined_branch_stall_in_signal))
			begin
				branch_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

module Matmul_basic_block_3
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_col_m2,
		input [63:0] 		input_rer,
		input [63:0] 		input_rei,
		input 		input_wii_cmp3,
		input 		valid_in,
		output 		stall_out,
		input 		input_exitcond,
		input [159:0] 		input_c0_exit_c0_exi4,
		input [31:0] 		input_c0_exe3,
		input [31:0] 		input_c0_exe4,
		input [31:0] 		input_global_id_0,
		input [31:0] 		input_global_id_1,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input 		start,
		input [255:0] 		avm_local_bb3_st_select40_readdata,
		input 		avm_local_bb3_st_select40_readdatavalid,
		input 		avm_local_bb3_st_select40_waitrequest,
		output [29:0] 		avm_local_bb3_st_select40_address,
		output 		avm_local_bb3_st_select40_read,
		output 		avm_local_bb3_st_select40_write,
		input 		avm_local_bb3_st_select40_writeack,
		output [255:0] 		avm_local_bb3_st_select40_writedata,
		output [31:0] 		avm_local_bb3_st_select40_byteenable,
		output [4:0] 		avm_local_bb3_st_select40_burstcount,
		output 		local_bb3_st_select40_active,
		input 		clock2x,
		input [255:0] 		avm_local_bb3_st_select37_readdata,
		input 		avm_local_bb3_st_select37_readdatavalid,
		input 		avm_local_bb3_st_select37_waitrequest,
		output [29:0] 		avm_local_bb3_st_select37_address,
		output 		avm_local_bb3_st_select37_read,
		output 		avm_local_bb3_st_select37_write,
		input 		avm_local_bb3_st_select37_writeack,
		output [255:0] 		avm_local_bb3_st_select37_writedata,
		output [31:0] 		avm_local_bb3_st_select37_byteenable,
		output [4:0] 		avm_local_bb3_st_select37_burstcount,
		output 		local_bb3_st_select37_active
	);


// Values used for debugging.  These are swept away by synthesis.
wire _entry;
wire _exit;
 reg [31:0] _num_entry_NO_SHIFT_REG;
 reg [31:0] _num_exit_NO_SHIFT_REG;
wire [31:0] _num_live;

assign _entry = ((&valid_in) & ~((|stall_out)));
assign _exit = ((&valid_out) & ~((|stall_in)));
assign _num_live = (_num_entry_NO_SHIFT_REG - _num_exit_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		_num_entry_NO_SHIFT_REG <= 32'h0;
		_num_exit_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		if (_entry)
		begin
			_num_entry_NO_SHIFT_REG <= (_num_entry_NO_SHIFT_REG + 2'h1);
		end
		if (_exit)
		begin
			_num_exit_NO_SHIFT_REG <= (_num_exit_NO_SHIFT_REG + 2'h1);
		end
	end
end



// This section defines the behaviour of the MERGE node
wire merge_node_stall_in_0;
 reg merge_node_valid_out_0_NO_SHIFT_REG;
wire merge_node_stall_in_1;
 reg merge_node_valid_out_1_NO_SHIFT_REG;
wire merge_node_stall_in_2;
 reg merge_node_valid_out_2_NO_SHIFT_REG;
wire merge_node_stall_in_3;
 reg merge_node_valid_out_3_NO_SHIFT_REG;
wire merge_node_stall_in_4;
 reg merge_node_valid_out_4_NO_SHIFT_REG;
wire merge_node_stall_in_5;
 reg merge_node_valid_out_5_NO_SHIFT_REG;
wire merge_stalled_by_successors;
 reg merge_block_selector_NO_SHIFT_REG;
 reg merge_node_valid_in_staging_reg_NO_SHIFT_REG;
 reg input_exitcond_staging_reg_NO_SHIFT_REG;
 reg [159:0] input_c0_exit_c0_exi4_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c0_exe3_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_c0_exe4_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_0_staging_reg_NO_SHIFT_REG;
 reg [31:0] input_global_id_1_staging_reg_NO_SHIFT_REG;
 reg local_lvm_exitcond_NO_SHIFT_REG;
 reg [159:0] local_lvm_c0_exit_c0_exi4_NO_SHIFT_REG;
 reg [31:0] local_lvm_c0_exe3_NO_SHIFT_REG;
 reg [31:0] local_lvm_c0_exe4_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_0_NO_SHIFT_REG;
 reg [31:0] local_lvm_input_global_id_1_NO_SHIFT_REG;
 reg is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
 reg invariant_valid_NO_SHIFT_REG;

assign merge_stalled_by_successors = ((merge_node_stall_in_0 & merge_node_valid_out_0_NO_SHIFT_REG) | (merge_node_stall_in_1 & merge_node_valid_out_1_NO_SHIFT_REG) | (merge_node_stall_in_2 & merge_node_valid_out_2_NO_SHIFT_REG) | (merge_node_stall_in_3 & merge_node_valid_out_3_NO_SHIFT_REG) | (merge_node_stall_in_4 & merge_node_valid_out_4_NO_SHIFT_REG) | (merge_node_stall_in_5 & merge_node_valid_out_5_NO_SHIFT_REG));
assign stall_out = merge_node_valid_in_staging_reg_NO_SHIFT_REG;

always @(*)
begin
	if ((merge_node_valid_in_staging_reg_NO_SHIFT_REG | valid_in))
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b1;
	end
	else
	begin
		merge_block_selector_NO_SHIFT_REG = 1'b0;
		is_merge_data_to_local_regs_valid_NO_SHIFT_REG = 1'b0;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		input_exitcond_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exit_c0_exi4_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe3_staging_reg_NO_SHIFT_REG <= 'x;
		input_c0_exe4_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_0_staging_reg_NO_SHIFT_REG <= 'x;
		input_global_id_1_staging_reg_NO_SHIFT_REG <= 'x;
		merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (((merge_block_selector_NO_SHIFT_REG != 1'b0) | merge_stalled_by_successors))
		begin
			if (~(merge_node_valid_in_staging_reg_NO_SHIFT_REG))
			begin
				input_exitcond_staging_reg_NO_SHIFT_REG <= input_exitcond;
				input_c0_exit_c0_exi4_staging_reg_NO_SHIFT_REG <= input_c0_exit_c0_exi4;
				input_c0_exe3_staging_reg_NO_SHIFT_REG <= input_c0_exe3;
				input_c0_exe4_staging_reg_NO_SHIFT_REG <= input_c0_exe4;
				input_global_id_0_staging_reg_NO_SHIFT_REG <= input_global_id_0;
				input_global_id_1_staging_reg_NO_SHIFT_REG <= input_global_id_1;
				merge_node_valid_in_staging_reg_NO_SHIFT_REG <= valid_in;
			end
		end
		else
		begin
			merge_node_valid_in_staging_reg_NO_SHIFT_REG <= 1'b0;
		end
	end
end

always @(posedge clock)
begin
	if (~(merge_stalled_by_successors))
	begin
		case (merge_block_selector_NO_SHIFT_REG)
			1'b0:
			begin
				if (merge_node_valid_in_staging_reg_NO_SHIFT_REG)
				begin
					local_lvm_exitcond_NO_SHIFT_REG <= input_exitcond_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exit_c0_exi4_NO_SHIFT_REG <= input_c0_exit_c0_exi4_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe3_NO_SHIFT_REG <= input_c0_exe3_staging_reg_NO_SHIFT_REG;
					local_lvm_c0_exe4_NO_SHIFT_REG <= input_c0_exe4_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0_staging_reg_NO_SHIFT_REG;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1_staging_reg_NO_SHIFT_REG;
				end
				else
				begin
					local_lvm_exitcond_NO_SHIFT_REG <= input_exitcond;
					local_lvm_c0_exit_c0_exi4_NO_SHIFT_REG <= input_c0_exit_c0_exi4;
					local_lvm_c0_exe3_NO_SHIFT_REG <= input_c0_exe3;
					local_lvm_c0_exe4_NO_SHIFT_REG <= input_c0_exe4;
					local_lvm_input_global_id_0_NO_SHIFT_REG <= input_global_id_0;
					local_lvm_input_global_id_1_NO_SHIFT_REG <= input_global_id_1;
				end
			end

			default:
			begin
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
		merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (~(merge_stalled_by_successors))
		begin
			merge_node_valid_out_0_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_1_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_2_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_3_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_4_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
			merge_node_valid_out_5_NO_SHIFT_REG <= is_merge_data_to_local_regs_valid_NO_SHIFT_REG;
		end
		else
		begin
			if (~(merge_node_stall_in_0))
			begin
				merge_node_valid_out_0_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_1))
			begin
				merge_node_valid_out_1_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_2))
			begin
				merge_node_valid_out_2_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_3))
			begin
				merge_node_valid_out_3_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_4))
			begin
				merge_node_valid_out_4_NO_SHIFT_REG <= 1'b0;
			end
			if (~(merge_node_stall_in_5))
			begin
				merge_node_valid_out_5_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		invariant_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		invariant_valid_NO_SHIFT_REG <= (~(start) & (invariant_valid_NO_SHIFT_REG | is_merge_data_to_local_regs_valid_NO_SHIFT_REG));
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe2_stall_local;
wire [31:0] local_bb3_c0_exe2;

assign local_bb3_c0_exe2 = local_lvm_c0_exit_c0_exi4_NO_SHIFT_REG[95:64];

// This section implements an unregistered operation.
// 
wire local_bb3_c0_exe1_stall_local;
wire [31:0] local_bb3_c0_exe1;

assign local_bb3_c0_exe1 = local_lvm_c0_exit_c0_exi4_NO_SHIFT_REG[63:32];

// This section implements a registered operation.
// 
wire local_bb3_mul40_inputs_ready;
 reg local_bb3_mul40_valid_out_NO_SHIFT_REG;
wire local_bb3_mul40_stall_in;
wire local_bb3_mul40_output_regs_ready;
wire [31:0] local_bb3_mul40;
 reg local_bb3_mul40_valid_pipe_0_NO_SHIFT_REG;
 reg local_bb3_mul40_valid_pipe_1_NO_SHIFT_REG;
wire local_bb3_mul40_causedstall;

acl_int_mult32s_s5 int_module_local_bb3_mul40 (
	.clock(clock),
	.dataa(local_lvm_input_global_id_1_NO_SHIFT_REG),
	.datab(input_col_m2),
	.enable(local_bb3_mul40_output_regs_ready),
	.result(local_bb3_mul40)
);

defparam int_module_local_bb3_mul40.INPUT1_WIDTH = 32;
defparam int_module_local_bb3_mul40.INPUT2_WIDTH = 32;

assign local_bb3_mul40_inputs_ready = merge_node_valid_out_4_NO_SHIFT_REG;
assign local_bb3_mul40_output_regs_ready = (&(~(local_bb3_mul40_valid_out_NO_SHIFT_REG) | ~(local_bb3_mul40_stall_in)));
assign merge_node_stall_in_4 = (~(local_bb3_mul40_output_regs_ready) | ~(local_bb3_mul40_inputs_ready));
assign local_bb3_mul40_causedstall = (local_bb3_mul40_inputs_ready && (~(local_bb3_mul40_output_regs_ready) && !(~(local_bb3_mul40_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul40_valid_pipe_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_mul40_valid_pipe_1_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul40_output_regs_ready)
		begin
			local_bb3_mul40_valid_pipe_0_NO_SHIFT_REG <= local_bb3_mul40_inputs_ready;
			local_bb3_mul40_valid_pipe_1_NO_SHIFT_REG <= local_bb3_mul40_valid_pipe_0_NO_SHIFT_REG;
		end
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_mul40_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_mul40_output_regs_ready)
		begin
			local_bb3_mul40_valid_out_NO_SHIFT_REG <= local_bb3_mul40_valid_pipe_1_NO_SHIFT_REG;
		end
		else
		begin
			if (~(local_bb3_mul40_stall_in))
			begin
				local_bb3_mul40_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// Register node:
//  * latency = 3
//  * capacity = 3
 logic rnode_1to4_input_global_id_0_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_1to4_input_global_id_0_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to4_input_global_id_0_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_1to4_input_global_id_0_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_lvm_input_global_id_0_NO_SHIFT_REG),
	.data_out(rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.DEPTH = 4;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to4_input_global_id_0_0_reg_4_fifo.IMPL = "ll_reg";

assign rnode_1to4_input_global_id_0_0_reg_4_inputs_ready_NO_SHIFT_REG = merge_node_valid_out_5_NO_SHIFT_REG;
assign merge_node_stall_in_5 = rnode_1to4_input_global_id_0_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_reg_4_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_stall_in_reg_4_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_stall_in_NO_SHIFT_REG;
assign rnode_1to4_input_global_id_0_0_valid_out_NO_SHIFT_REG = rnode_1to4_input_global_id_0_0_valid_out_reg_4_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__31_stall_local;
wire [31:0] local_bb3__31;

assign local_bb3__31 = (local_lvm_exitcond_NO_SHIFT_REG ? local_bb3_c0_exe2 : local_lvm_c0_exe4_NO_SHIFT_REG);

// This section implements an unregistered operation.
// 
wire local_bb3__33_stall_local;
wire [31:0] local_bb3__33;

assign local_bb3__33 = (local_lvm_exitcond_NO_SHIFT_REG ? local_bb3_c0_exe1 : local_lvm_c0_exe3_NO_SHIFT_REG);

// Register node:
//  * latency = 0
//  * capacity = 2
 logic rnode_4to4_bb3_mul40_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to4_bb3_mul40_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb3_mul40_0_NO_SHIFT_REG;
 logic rnode_4to4_bb3_mul40_0_reg_4_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to4_bb3_mul40_0_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb3_mul40_0_valid_out_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb3_mul40_0_stall_in_reg_4_NO_SHIFT_REG;
 logic rnode_4to4_bb3_mul40_0_stall_out_reg_4_NO_SHIFT_REG;

acl_data_fifo rnode_4to4_bb3_mul40_0_reg_4_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to4_bb3_mul40_0_reg_4_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to4_bb3_mul40_0_stall_in_reg_4_NO_SHIFT_REG),
	.valid_out(rnode_4to4_bb3_mul40_0_valid_out_reg_4_NO_SHIFT_REG),
	.stall_out(rnode_4to4_bb3_mul40_0_stall_out_reg_4_NO_SHIFT_REG),
	.data_in(local_bb3_mul40),
	.data_out(rnode_4to4_bb3_mul40_0_reg_4_NO_SHIFT_REG)
);

defparam rnode_4to4_bb3_mul40_0_reg_4_fifo.DEPTH = 3;
defparam rnode_4to4_bb3_mul40_0_reg_4_fifo.DATA_WIDTH = 32;
defparam rnode_4to4_bb3_mul40_0_reg_4_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to4_bb3_mul40_0_reg_4_fifo.IMPL = "zl_reg";

assign rnode_4to4_bb3_mul40_0_reg_4_inputs_ready_NO_SHIFT_REG = local_bb3_mul40_valid_out_NO_SHIFT_REG;
assign local_bb3_mul40_stall_in = rnode_4to4_bb3_mul40_0_stall_out_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb3_mul40_0_NO_SHIFT_REG = rnode_4to4_bb3_mul40_0_reg_4_NO_SHIFT_REG;
assign rnode_4to4_bb3_mul40_0_stall_in_reg_4_NO_SHIFT_REG = rnode_4to4_bb3_mul40_0_stall_in_NO_SHIFT_REG;
assign rnode_4to4_bb3_mul40_0_valid_out_NO_SHIFT_REG = rnode_4to4_bb3_mul40_0_valid_out_reg_4_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_var__stall_local;
wire [31:0] local_bb3_var_;

assign local_bb3_var_ = local_bb3__31;

// This section implements an unregistered operation.
// 
wire local_bb3_var__u176_stall_local;
wire [31:0] local_bb3_var__u176;

assign local_bb3_var__u176 = local_bb3__33;

// This section implements an unregistered operation.
// 
wire local_bb3_add41_valid_out;
wire local_bb3_add41_stall_in;
wire local_bb3_add41_inputs_ready;
wire local_bb3_add41_stall_local;
wire [31:0] local_bb3_add41;

assign local_bb3_add41_inputs_ready = (rnode_1to4_input_global_id_0_0_valid_out_NO_SHIFT_REG & rnode_4to4_bb3_mul40_0_valid_out_NO_SHIFT_REG);
assign local_bb3_add41 = (rnode_4to4_bb3_mul40_0_NO_SHIFT_REG + rnode_1to4_input_global_id_0_0_NO_SHIFT_REG);
assign local_bb3_add41_valid_out = local_bb3_add41_inputs_ready;
assign local_bb3_add41_stall_local = local_bb3_add41_stall_in;
assign rnode_1to4_input_global_id_0_0_stall_in_NO_SHIFT_REG = (local_bb3_add41_stall_local | ~(local_bb3_add41_inputs_ready));
assign rnode_4to4_bb3_mul40_0_stall_in_NO_SHIFT_REG = (local_bb3_add41_stall_local | ~(local_bb3_add41_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i1_stall_local;
wire [31:0] local_bb3_shr_i1;

assign local_bb3_shr_i1 = (local_bb3_var_ >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and2_i_stall_local;
wire [31:0] local_bb3_and2_i;

assign local_bb3_and2_i = (local_bb3_var_ & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and33_i_stall_local;
wire [31:0] local_bb3_and33_i;

assign local_bb3_and33_i = (local_bb3_var_ & 32'h807FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_shr_i7_stall_local;
wire [31:0] local_bb3_shr_i7;

assign local_bb3_shr_i7 = (local_bb3_var__u176 >> 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_and2_i10_stall_local;
wire [31:0] local_bb3_and2_i10;

assign local_bb3_and2_i10 = (local_bb3_var__u176 & 32'h7FFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_and33_i34_stall_local;
wire [31:0] local_bb3_and33_i34;

assign local_bb3_and33_i34 = (local_bb3_var__u176 & 32'h807FFFFF);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_4to5_bb3_add41_0_valid_out_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add41_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_add41_0_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add41_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_4to5_bb3_add41_0_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add41_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add41_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_4to5_bb3_add41_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_4to5_bb3_add41_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_4to5_bb3_add41_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_4to5_bb3_add41_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_4to5_bb3_add41_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_4to5_bb3_add41_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_add41),
	.data_out(rnode_4to5_bb3_add41_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_4to5_bb3_add41_0_reg_5_fifo.DEPTH = 2;
defparam rnode_4to5_bb3_add41_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_4to5_bb3_add41_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_4to5_bb3_add41_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_4to5_bb3_add41_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb3_add41_valid_out;
assign local_bb3_add41_stall_in = rnode_4to5_bb3_add41_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_add41_0_NO_SHIFT_REG = rnode_4to5_bb3_add41_0_reg_5_NO_SHIFT_REG;
assign rnode_4to5_bb3_add41_0_stall_in_reg_5_NO_SHIFT_REG = rnode_4to5_bb3_add41_0_stall_in_NO_SHIFT_REG;
assign rnode_4to5_bb3_add41_0_valid_out_NO_SHIFT_REG = rnode_4to5_bb3_add41_0_valid_out_reg_5_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_and1_i_stall_local;
wire [31:0] local_bb3_and1_i;

assign local_bb3_and1_i = (local_bb3_shr_i1 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot6_i_stall_local;
wire local_bb3_lnot6_i;

assign local_bb3_lnot6_i = (local_bb3_and2_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and1_i8_stall_local;
wire [31:0] local_bb3_and1_i8;

assign local_bb3_and1_i8 = (local_bb3_shr_i7 & 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_lnot6_i11_stall_local;
wire local_bb3_lnot6_i11;

assign local_bb3_lnot6_i11 = (local_bb3_and2_i10 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_idxprom42_stall_local;
wire [63:0] local_bb3_idxprom42;

assign local_bb3_idxprom42[32] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[33] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[34] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[35] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[36] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[37] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[38] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[39] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[40] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[41] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[42] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[43] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[44] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[45] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[46] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[47] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[48] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[49] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[50] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[51] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[52] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[53] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[54] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[55] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[56] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[57] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[58] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[59] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[60] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[61] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[62] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[63] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG[31];
assign local_bb3_idxprom42[31:0] = rnode_4to5_bb3_add41_0_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i2_stall_local;
wire local_bb3_cmp_i2;

assign local_bb3_cmp_i2 = (local_bb3_and1_i == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp10_i_stall_local;
wire local_bb3_cmp10_i;

assign local_bb3_cmp10_i = (local_bb3_and1_i == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp_i9_stall_local;
wire local_bb3_cmp_i9;

assign local_bb3_cmp_i9 = (local_bb3_and1_i8 == 32'hFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp10_i12_stall_local;
wire local_bb3_cmp10_i12;

assign local_bb3_cmp10_i12 = (local_bb3_and1_i8 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_arrayidx43_stall_local;
wire [63:0] local_bb3_arrayidx43;

assign local_bb3_arrayidx43 = (input_rer + (local_bb3_idxprom42 << 6'h2));

// This section implements an unregistered operation.
// 
wire local_bb3_arrayidx43_valid_out;
wire local_bb3_arrayidx43_stall_in;
 reg local_bb3_arrayidx43_consumed_0_NO_SHIFT_REG;
wire local_bb3_arrayidx48_valid_out;
wire local_bb3_arrayidx48_stall_in;
 reg local_bb3_arrayidx48_consumed_0_NO_SHIFT_REG;
wire local_bb3_arrayidx48_inputs_ready;
wire local_bb3_arrayidx48_stall_local;
wire [63:0] local_bb3_arrayidx48;

assign local_bb3_arrayidx48_inputs_ready = rnode_4to5_bb3_add41_0_valid_out_NO_SHIFT_REG;
assign local_bb3_arrayidx48 = (input_rei + (local_bb3_idxprom42 << 6'h2));
assign local_bb3_arrayidx48_stall_local = ((local_bb3_arrayidx43_stall_in & ~(local_bb3_arrayidx43_consumed_0_NO_SHIFT_REG)) | (local_bb3_arrayidx48_stall_in & ~(local_bb3_arrayidx48_consumed_0_NO_SHIFT_REG)));
assign local_bb3_arrayidx43_valid_out = (local_bb3_arrayidx48_inputs_ready & ~(local_bb3_arrayidx43_consumed_0_NO_SHIFT_REG));
assign local_bb3_arrayidx48_valid_out = (local_bb3_arrayidx48_inputs_ready & ~(local_bb3_arrayidx48_consumed_0_NO_SHIFT_REG));
assign rnode_4to5_bb3_add41_0_stall_in_NO_SHIFT_REG = (|local_bb3_arrayidx48_stall_local);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_arrayidx43_consumed_0_NO_SHIFT_REG <= 1'b0;
		local_bb3_arrayidx48_consumed_0_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		local_bb3_arrayidx43_consumed_0_NO_SHIFT_REG <= (local_bb3_arrayidx48_inputs_ready & (local_bb3_arrayidx43_consumed_0_NO_SHIFT_REG | ~(local_bb3_arrayidx43_stall_in)) & local_bb3_arrayidx48_stall_local);
		local_bb3_arrayidx48_consumed_0_NO_SHIFT_REG <= (local_bb3_arrayidx48_inputs_ready & (local_bb3_arrayidx48_consumed_0_NO_SHIFT_REG | ~(local_bb3_arrayidx48_stall_in)) & local_bb3_arrayidx48_stall_local);
	end
end


// This section implements an unregistered operation.
// 
wire local_bb3___i_stall_local;
wire local_bb3___i;

assign local_bb3___i = (local_bb3_cmp_i2 & local_bb3_lnot6_i);

// This section implements an unregistered operation.
// 
wire local_bb3_not_cmp_i_stall_local;
wire local_bb3_not_cmp_i;

assign local_bb3_not_cmp_i = (local_bb3_cmp_i2 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_conv22_i_stall_local;
wire [31:0] local_bb3_conv22_i;

assign local_bb3_conv22_i[31:1] = 31'h0;
assign local_bb3_conv22_i[0] = local_bb3_cmp_i2;

// This section implements an unregistered operation.
// 
wire local_bb3_not_cmp10_i_stall_local;
wire local_bb3_not_cmp10_i;

assign local_bb3_not_cmp10_i = (local_bb3_cmp10_i ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3___i13_stall_local;
wire local_bb3___i13;

assign local_bb3___i13 = (local_bb3_cmp_i9 & local_bb3_lnot6_i11);

// This section implements an unregistered operation.
// 
wire local_bb3_not_cmp_i14_stall_local;
wire local_bb3_not_cmp_i14;

assign local_bb3_not_cmp_i14 = (local_bb3_cmp_i9 ^ 1'b1);

// This section implements an unregistered operation.
// 
wire local_bb3_conv22_i29_stall_local;
wire [31:0] local_bb3_conv22_i29;

assign local_bb3_conv22_i29[31:1] = 31'h0;
assign local_bb3_conv22_i29[0] = local_bb3_cmp_i9;

// This section implements an unregistered operation.
// 
wire local_bb3_not_cmp10_i17_stall_local;
wire local_bb3_not_cmp10_i17;

assign local_bb3_not_cmp10_i17 = (local_bb3_cmp10_i12 ^ 1'b1);

// This section implements a staging register.
// 
wire rstag_5to5_bb3_arrayidx43_valid_out;
wire rstag_5to5_bb3_arrayidx43_stall_in;
wire rstag_5to5_bb3_arrayidx43_inputs_ready;
wire rstag_5to5_bb3_arrayidx43_stall_local;
 reg rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG;
wire rstag_5to5_bb3_arrayidx43_combined_valid;
 reg [63:0] rstag_5to5_bb3_arrayidx43_staging_reg_NO_SHIFT_REG;
wire [63:0] rstag_5to5_bb3_arrayidx43;

assign rstag_5to5_bb3_arrayidx43_inputs_ready = local_bb3_arrayidx43_valid_out;
assign rstag_5to5_bb3_arrayidx43 = (rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG ? rstag_5to5_bb3_arrayidx43_staging_reg_NO_SHIFT_REG : local_bb3_arrayidx43);
assign rstag_5to5_bb3_arrayidx43_combined_valid = (rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG | rstag_5to5_bb3_arrayidx43_inputs_ready);
assign rstag_5to5_bb3_arrayidx43_valid_out = rstag_5to5_bb3_arrayidx43_combined_valid;
assign rstag_5to5_bb3_arrayidx43_stall_local = rstag_5to5_bb3_arrayidx43_stall_in;
assign local_bb3_arrayidx43_stall_in = (|rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_5to5_bb3_arrayidx43_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_5to5_bb3_arrayidx43_stall_local)
		begin
			if (~(rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG))
			begin
				rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG <= rstag_5to5_bb3_arrayidx43_inputs_ready;
			end
		end
		else
		begin
			rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_5to5_bb3_arrayidx43_staging_valid_NO_SHIFT_REG))
		begin
			rstag_5to5_bb3_arrayidx43_staging_reg_NO_SHIFT_REG <= local_bb3_arrayidx43;
		end
	end
end


// Register node:
//  * latency = 137
//  * capacity = 137
 logic rnode_5to142_bb3_arrayidx48_0_valid_out_NO_SHIFT_REG;
 logic rnode_5to142_bb3_arrayidx48_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_5to142_bb3_arrayidx48_0_NO_SHIFT_REG;
 logic rnode_5to142_bb3_arrayidx48_0_reg_142_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_5to142_bb3_arrayidx48_0_reg_142_NO_SHIFT_REG;
 logic rnode_5to142_bb3_arrayidx48_0_valid_out_reg_142_NO_SHIFT_REG;
 logic rnode_5to142_bb3_arrayidx48_0_stall_in_reg_142_NO_SHIFT_REG;
 logic rnode_5to142_bb3_arrayidx48_0_stall_out_reg_142_NO_SHIFT_REG;

acl_data_fifo rnode_5to142_bb3_arrayidx48_0_reg_142_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_5to142_bb3_arrayidx48_0_reg_142_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_5to142_bb3_arrayidx48_0_stall_in_reg_142_NO_SHIFT_REG),
	.valid_out(rnode_5to142_bb3_arrayidx48_0_valid_out_reg_142_NO_SHIFT_REG),
	.stall_out(rnode_5to142_bb3_arrayidx48_0_stall_out_reg_142_NO_SHIFT_REG),
	.data_in(local_bb3_arrayidx48),
	.data_out(rnode_5to142_bb3_arrayidx48_0_reg_142_NO_SHIFT_REG)
);

defparam rnode_5to142_bb3_arrayidx48_0_reg_142_fifo.DEPTH = 138;
defparam rnode_5to142_bb3_arrayidx48_0_reg_142_fifo.DATA_WIDTH = 64;
defparam rnode_5to142_bb3_arrayidx48_0_reg_142_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_5to142_bb3_arrayidx48_0_reg_142_fifo.IMPL = "ram";

assign rnode_5to142_bb3_arrayidx48_0_reg_142_inputs_ready_NO_SHIFT_REG = local_bb3_arrayidx48_valid_out;
assign local_bb3_arrayidx48_stall_in = rnode_5to142_bb3_arrayidx48_0_stall_out_reg_142_NO_SHIFT_REG;
assign rnode_5to142_bb3_arrayidx48_0_NO_SHIFT_REG = rnode_5to142_bb3_arrayidx48_0_reg_142_NO_SHIFT_REG;
assign rnode_5to142_bb3_arrayidx48_0_stall_in_reg_142_NO_SHIFT_REG = rnode_5to142_bb3_arrayidx48_0_stall_in_NO_SHIFT_REG;
assign rnode_5to142_bb3_arrayidx48_0_valid_out_NO_SHIFT_REG = rnode_5to142_bb3_arrayidx48_0_valid_out_reg_142_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_conv44_i_stall_local;
wire [31:0] local_bb3_conv44_i;

assign local_bb3_conv44_i[31:1] = 31'h0;
assign local_bb3_conv44_i[0] = local_bb3___i;

// This section implements an unregistered operation.
// 
wire local_bb3_cond50_i_stall_local;
wire [31:0] local_bb3_cond50_i;

assign local_bb3_cond50_i = (local_bb3___i ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__4_i_stall_local;
wire local_bb3__4_i;

assign local_bb3__4_i = (local_bb3_cmp10_i & local_bb3_not_cmp_i);

// This section implements an unregistered operation.
// 
wire local_bb3__7_i_stall_local;
wire local_bb3__7_i;

assign local_bb3__7_i = (local_bb3_cmp_i2 | local_bb3_not_cmp10_i);

// This section implements an unregistered operation.
// 
wire local_bb3_conv44_i42_stall_local;
wire [31:0] local_bb3_conv44_i42;

assign local_bb3_conv44_i42[31:1] = 31'h0;
assign local_bb3_conv44_i42[0] = local_bb3___i13;

// This section implements an unregistered operation.
// 
wire local_bb3_cond50_i46_stall_local;
wire [31:0] local_bb3_cond50_i46;

assign local_bb3_cond50_i46 = (local_bb3___i13 ? 32'h400000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3__4_i15_stall_local;
wire local_bb3__4_i15;

assign local_bb3__4_i15 = (local_bb3_cmp10_i12 & local_bb3_not_cmp_i14);

// This section implements an unregistered operation.
// 
wire local_bb3__7_i18_stall_local;
wire local_bb3__7_i18;

assign local_bb3__7_i18 = (local_bb3_cmp_i9 | local_bb3_not_cmp10_i17);

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_142to143_bb3_arrayidx48_0_valid_out_NO_SHIFT_REG;
 logic rnode_142to143_bb3_arrayidx48_0_stall_in_NO_SHIFT_REG;
 logic [63:0] rnode_142to143_bb3_arrayidx48_0_NO_SHIFT_REG;
 logic rnode_142to143_bb3_arrayidx48_0_reg_143_inputs_ready_NO_SHIFT_REG;
 logic [63:0] rnode_142to143_bb3_arrayidx48_0_reg_143_NO_SHIFT_REG;
 logic rnode_142to143_bb3_arrayidx48_0_valid_out_reg_143_NO_SHIFT_REG;
 logic rnode_142to143_bb3_arrayidx48_0_stall_in_reg_143_NO_SHIFT_REG;
 logic rnode_142to143_bb3_arrayidx48_0_stall_out_reg_143_NO_SHIFT_REG;

acl_data_fifo rnode_142to143_bb3_arrayidx48_0_reg_143_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_142to143_bb3_arrayidx48_0_reg_143_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_142to143_bb3_arrayidx48_0_stall_in_reg_143_NO_SHIFT_REG),
	.valid_out(rnode_142to143_bb3_arrayidx48_0_valid_out_reg_143_NO_SHIFT_REG),
	.stall_out(rnode_142to143_bb3_arrayidx48_0_stall_out_reg_143_NO_SHIFT_REG),
	.data_in(rnode_5to142_bb3_arrayidx48_0_NO_SHIFT_REG),
	.data_out(rnode_142to143_bb3_arrayidx48_0_reg_143_NO_SHIFT_REG)
);

defparam rnode_142to143_bb3_arrayidx48_0_reg_143_fifo.DEPTH = 2;
defparam rnode_142to143_bb3_arrayidx48_0_reg_143_fifo.DATA_WIDTH = 64;
defparam rnode_142to143_bb3_arrayidx48_0_reg_143_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_142to143_bb3_arrayidx48_0_reg_143_fifo.IMPL = "ll_reg";

assign rnode_142to143_bb3_arrayidx48_0_reg_143_inputs_ready_NO_SHIFT_REG = rnode_5to142_bb3_arrayidx48_0_valid_out_NO_SHIFT_REG;
assign rnode_5to142_bb3_arrayidx48_0_stall_in_NO_SHIFT_REG = rnode_142to143_bb3_arrayidx48_0_stall_out_reg_143_NO_SHIFT_REG;
assign rnode_142to143_bb3_arrayidx48_0_NO_SHIFT_REG = rnode_142to143_bb3_arrayidx48_0_reg_143_NO_SHIFT_REG;
assign rnode_142to143_bb3_arrayidx48_0_stall_in_reg_143_NO_SHIFT_REG = rnode_142to143_bb3_arrayidx48_0_stall_in_NO_SHIFT_REG;
assign rnode_142to143_bb3_arrayidx48_0_valid_out_NO_SHIFT_REG = rnode_142to143_bb3_arrayidx48_0_valid_out_reg_143_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3__5_i_stall_local;
wire [31:0] local_bb3__5_i;

assign local_bb3__5_i[31:1] = 31'h0;
assign local_bb3__5_i[0] = local_bb3__4_i;

// This section implements an unregistered operation.
// 
wire local_bb3__17_i_stall_local;
wire [31:0] local_bb3__17_i;

assign local_bb3__17_i = (local_bb3__4_i ? 32'h0 : 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb3__5_i16_stall_local;
wire [31:0] local_bb3__5_i16;

assign local_bb3__5_i16[31:1] = 31'h0;
assign local_bb3__5_i16[0] = local_bb3__4_i15;

// This section implements an unregistered operation.
// 
wire local_bb3__17_i23_stall_local;
wire [31:0] local_bb3__17_i23;

assign local_bb3__17_i23 = (local_bb3__4_i15 ? 32'h0 : 32'h100);

// This section implements an unregistered operation.
// 
wire local_bb3__9_i_stall_local;
wire [31:0] local_bb3__9_i;

assign local_bb3__9_i = (local_bb3__7_i ? 32'h0 : local_bb3__5_i);

// This section implements an unregistered operation.
// 
wire local_bb3__18_i_stall_local;
wire [31:0] local_bb3__18_i;

assign local_bb3__18_i = (local_bb3__7_i ? 32'h0 : local_bb3__17_i);

// This section implements an unregistered operation.
// 
wire local_bb3__9_i20_stall_local;
wire [31:0] local_bb3__9_i20;

assign local_bb3__9_i20 = (local_bb3__7_i18 ? 32'h0 : local_bb3__5_i16);

// This section implements an unregistered operation.
// 
wire local_bb3__18_i24_stall_local;
wire [31:0] local_bb3__18_i24;

assign local_bb3__18_i24 = (local_bb3__7_i18 ? 32'h0 : local_bb3__17_i23);

// This section implements an unregistered operation.
// 
wire local_bb3_add_i3_stall_local;
wire [31:0] local_bb3_add_i3;

assign local_bb3_add_i3 = (local_bb3__18_i | local_bb3_and1_i);

// This section implements an unregistered operation.
// 
wire local_bb3_fold_i_stall_local;
wire [31:0] local_bb3_fold_i;

assign local_bb3_fold_i = (local_bb3__18_i + local_bb3_shr_i1);

// This section implements an unregistered operation.
// 
wire local_bb3_add_i26_stall_local;
wire [31:0] local_bb3_add_i26;

assign local_bb3_add_i26 = (local_bb3__18_i24 | local_bb3_and1_i8);

// This section implements an unregistered operation.
// 
wire local_bb3_fold_i33_stall_local;
wire [31:0] local_bb3_fold_i33;

assign local_bb3_fold_i33 = (local_bb3__18_i24 + local_bb3_shr_i7);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp20_i_stall_local;
wire local_bb3_cmp20_i;

assign local_bb3_cmp20_i = (local_bb3_add_i3 > 32'hFE);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp25_i_stall_local;
wire local_bb3_cmp25_i;

assign local_bb3_cmp25_i = (local_bb3_add_i3 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and32_i_stall_local;
wire [31:0] local_bb3_and32_i;

assign local_bb3_and32_i = (local_bb3_fold_i << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp20_i27_stall_local;
wire local_bb3_cmp20_i27;

assign local_bb3_cmp20_i27 = (local_bb3_add_i26 > 32'hFE);

// This section implements an unregistered operation.
// 
wire local_bb3_cmp25_i31_stall_local;
wire local_bb3_cmp25_i31;

assign local_bb3_cmp25_i31 = (local_bb3_add_i26 == 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_and32_i35_stall_local;
wire [31:0] local_bb3_and32_i35;

assign local_bb3_and32_i35 = (local_bb3_fold_i33 << 32'h17);

// This section implements an unregistered operation.
// 
wire local_bb3_conv_i_stall_local;
wire [31:0] local_bb3_conv_i;

assign local_bb3_conv_i[31:1] = 31'h0;
assign local_bb3_conv_i[0] = local_bb3_cmp20_i;

// This section implements an unregistered operation.
// 
wire local_bb3_conv26_i_stall_local;
wire [31:0] local_bb3_conv26_i;

assign local_bb3_conv26_i[31:1] = 31'h0;
assign local_bb3_conv26_i[0] = local_bb3_cmp25_i;

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i5_stall_local;
wire [31:0] local_bb3_shl_i5;

assign local_bb3_shl_i5 = (local_bb3_and32_i & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb3_conv_i28_stall_local;
wire [31:0] local_bb3_conv_i28;

assign local_bb3_conv_i28[31:1] = 31'h0;
assign local_bb3_conv_i28[0] = local_bb3_cmp20_i27;

// This section implements an unregistered operation.
// 
wire local_bb3_conv26_i32_stall_local;
wire [31:0] local_bb3_conv26_i32;

assign local_bb3_conv26_i32[31:1] = 31'h0;
assign local_bb3_conv26_i32[0] = local_bb3_cmp25_i31;

// This section implements an unregistered operation.
// 
wire local_bb3_shl_i36_stall_local;
wire [31:0] local_bb3_shl_i36;

assign local_bb3_shl_i36 = (local_bb3_and32_i35 & 32'h7F800000);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i4_stall_local;
wire [31:0] local_bb3_or_i4;

assign local_bb3_or_i4 = (local_bb3_conv_i | local_bb3_conv22_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or29_i_stall_local;
wire [31:0] local_bb3_or29_i;

assign local_bb3_or29_i = (local_bb3_conv26_i | local_bb3__9_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or34_i_stall_local;
wire [31:0] local_bb3_or34_i;

assign local_bb3_or34_i = (local_bb3_shl_i5 | local_bb3_and33_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or_i30_stall_local;
wire [31:0] local_bb3_or_i30;

assign local_bb3_or_i30 = (local_bb3_conv_i28 | local_bb3_conv22_i29);

// This section implements an unregistered operation.
// 
wire local_bb3_or29_i38_stall_local;
wire [31:0] local_bb3_or29_i38;

assign local_bb3_or29_i38 = (local_bb3_conv26_i32 | local_bb3__9_i20);

// This section implements an unregistered operation.
// 
wire local_bb3_or34_i37_stall_local;
wire [31:0] local_bb3_or34_i37;

assign local_bb3_or34_i37 = (local_bb3_shl_i36 | local_bb3_and33_i34);

// This section implements an unregistered operation.
// 
wire local_bb3_or45_i_stall_local;
wire [31:0] local_bb3_or45_i;

assign local_bb3_or45_i = (local_bb3_or_i4 | local_bb3_conv44_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or39_i_stall_local;
wire [31:0] local_bb3_or39_i;

assign local_bb3_or39_i = (local_bb3_or29_i | local_bb3_or_i4);

// This section implements an unregistered operation.
// 
wire local_bb3_or45_i43_stall_local;
wire [31:0] local_bb3_or45_i43;

assign local_bb3_or45_i43 = (local_bb3_or_i30 | local_bb3_conv44_i42);

// This section implements an unregistered operation.
// 
wire local_bb3_or39_i39_stall_local;
wire [31:0] local_bb3_or39_i39;

assign local_bb3_or39_i39 = (local_bb3_or29_i38 | local_bb3_or_i30);

// This section implements an unregistered operation.
// 
wire local_bb3_tobool46_i_stall_local;
wire local_bb3_tobool46_i;

assign local_bb3_tobool46_i = (local_bb3_or45_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_tobool40_i_stall_local;
wire local_bb3_tobool40_i;

assign local_bb3_tobool40_i = (local_bb3_or39_i != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_tobool46_i44_stall_local;
wire local_bb3_tobool46_i44;

assign local_bb3_tobool46_i44 = (local_bb3_or45_i43 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_tobool40_i40_stall_local;
wire local_bb3_tobool40_i40;

assign local_bb3_tobool40_i40 = (local_bb3_or39_i39 != 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cond47_i_stall_local;
wire [31:0] local_bb3_cond47_i;

assign local_bb3_cond47_i = (local_bb3_tobool46_i ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cond_i6_stall_local;
wire [31:0] local_bb3_cond_i6;

assign local_bb3_cond_i6 = (local_bb3_tobool40_i ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_cond47_i45_stall_local;
wire [31:0] local_bb3_cond47_i45;

assign local_bb3_cond47_i45 = (local_bb3_tobool46_i44 ? 32'h7F800000 : 32'h0);

// This section implements an unregistered operation.
// 
wire local_bb3_cond_i41_stall_local;
wire [31:0] local_bb3_cond_i41;

assign local_bb3_cond_i41 = (local_bb3_tobool40_i40 ? 32'h80000000 : 32'hFFFFFFFF);

// This section implements an unregistered operation.
// 
wire local_bb3_or52_i_stall_local;
wire [31:0] local_bb3_or52_i;

assign local_bb3_or52_i = (local_bb3_cond47_i | local_bb3_cond50_i);

// This section implements an unregistered operation.
// 
wire local_bb3_and51_i_stall_local;
wire [31:0] local_bb3_and51_i;

assign local_bb3_and51_i = (local_bb3_cond_i6 & local_bb3_or34_i);

// This section implements an unregistered operation.
// 
wire local_bb3_or52_i48_stall_local;
wire [31:0] local_bb3_or52_i48;

assign local_bb3_or52_i48 = (local_bb3_cond47_i45 | local_bb3_cond50_i46);

// This section implements an unregistered operation.
// 
wire local_bb3_and51_i47_stall_local;
wire [31:0] local_bb3_and51_i47;

assign local_bb3_and51_i47 = (local_bb3_cond_i41 & local_bb3_or34_i37);

// This section implements an unregistered operation.
// 
wire local_bb3_or53_i_valid_out;
wire local_bb3_or53_i_stall_in;
wire local_bb3_or53_i_inputs_ready;
wire local_bb3_or53_i_stall_local;
wire [31:0] local_bb3_or53_i;

assign local_bb3_or53_i_inputs_ready = (merge_node_valid_out_0_NO_SHIFT_REG & merge_node_valid_out_2_NO_SHIFT_REG);
assign local_bb3_or53_i = (local_bb3_or52_i | local_bb3_and51_i);
assign local_bb3_or53_i_valid_out = local_bb3_or53_i_inputs_ready;
assign local_bb3_or53_i_stall_local = local_bb3_or53_i_stall_in;
assign merge_node_stall_in_0 = (local_bb3_or53_i_stall_local | ~(local_bb3_or53_i_inputs_ready));
assign merge_node_stall_in_2 = (local_bb3_or53_i_stall_local | ~(local_bb3_or53_i_inputs_ready));

// This section implements an unregistered operation.
// 
wire local_bb3_or53_i49_valid_out;
wire local_bb3_or53_i49_stall_in;
wire local_bb3_or53_i49_inputs_ready;
wire local_bb3_or53_i49_stall_local;
wire [31:0] local_bb3_or53_i49;

assign local_bb3_or53_i49_inputs_ready = (merge_node_valid_out_1_NO_SHIFT_REG & merge_node_valid_out_3_NO_SHIFT_REG);
assign local_bb3_or53_i49 = (local_bb3_or52_i48 | local_bb3_and51_i47);
assign local_bb3_or53_i49_valid_out = local_bb3_or53_i49_inputs_ready;
assign local_bb3_or53_i49_stall_local = local_bb3_or53_i49_stall_in;
assign merge_node_stall_in_1 = (local_bb3_or53_i49_stall_local | ~(local_bb3_or53_i49_inputs_ready));
assign merge_node_stall_in_3 = (local_bb3_or53_i49_stall_local | ~(local_bb3_or53_i49_inputs_ready));

// Register node:
//  * latency = 141
//  * capacity = 141
 logic rnode_1to142_bb3_or53_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to142_bb3_or53_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to142_bb3_or53_i_0_NO_SHIFT_REG;
 logic rnode_1to142_bb3_or53_i_0_reg_142_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to142_bb3_or53_i_0_reg_142_NO_SHIFT_REG;
 logic rnode_1to142_bb3_or53_i_0_valid_out_reg_142_NO_SHIFT_REG;
 logic rnode_1to142_bb3_or53_i_0_stall_in_reg_142_NO_SHIFT_REG;
 logic rnode_1to142_bb3_or53_i_0_stall_out_reg_142_NO_SHIFT_REG;

acl_data_fifo rnode_1to142_bb3_or53_i_0_reg_142_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to142_bb3_or53_i_0_reg_142_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to142_bb3_or53_i_0_stall_in_reg_142_NO_SHIFT_REG),
	.valid_out(rnode_1to142_bb3_or53_i_0_valid_out_reg_142_NO_SHIFT_REG),
	.stall_out(rnode_1to142_bb3_or53_i_0_stall_out_reg_142_NO_SHIFT_REG),
	.data_in(local_bb3_or53_i),
	.data_out(rnode_1to142_bb3_or53_i_0_reg_142_NO_SHIFT_REG)
);

defparam rnode_1to142_bb3_or53_i_0_reg_142_fifo.DEPTH = 142;
defparam rnode_1to142_bb3_or53_i_0_reg_142_fifo.DATA_WIDTH = 32;
defparam rnode_1to142_bb3_or53_i_0_reg_142_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to142_bb3_or53_i_0_reg_142_fifo.IMPL = "ram";

assign rnode_1to142_bb3_or53_i_0_reg_142_inputs_ready_NO_SHIFT_REG = local_bb3_or53_i_valid_out;
assign local_bb3_or53_i_stall_in = rnode_1to142_bb3_or53_i_0_stall_out_reg_142_NO_SHIFT_REG;
assign rnode_1to142_bb3_or53_i_0_NO_SHIFT_REG = rnode_1to142_bb3_or53_i_0_reg_142_NO_SHIFT_REG;
assign rnode_1to142_bb3_or53_i_0_stall_in_reg_142_NO_SHIFT_REG = rnode_1to142_bb3_or53_i_0_stall_in_NO_SHIFT_REG;
assign rnode_1to142_bb3_or53_i_0_valid_out_NO_SHIFT_REG = rnode_1to142_bb3_or53_i_0_valid_out_reg_142_NO_SHIFT_REG;

// Register node:
//  * latency = 4
//  * capacity = 4
 logic rnode_1to5_bb3_or53_i49_0_valid_out_NO_SHIFT_REG;
 logic rnode_1to5_bb3_or53_i49_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_1to5_bb3_or53_i49_0_NO_SHIFT_REG;
 logic rnode_1to5_bb3_or53_i49_0_reg_5_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_1to5_bb3_or53_i49_0_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb3_or53_i49_0_valid_out_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb3_or53_i49_0_stall_in_reg_5_NO_SHIFT_REG;
 logic rnode_1to5_bb3_or53_i49_0_stall_out_reg_5_NO_SHIFT_REG;

acl_data_fifo rnode_1to5_bb3_or53_i49_0_reg_5_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_1to5_bb3_or53_i49_0_reg_5_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_1to5_bb3_or53_i49_0_stall_in_reg_5_NO_SHIFT_REG),
	.valid_out(rnode_1to5_bb3_or53_i49_0_valid_out_reg_5_NO_SHIFT_REG),
	.stall_out(rnode_1to5_bb3_or53_i49_0_stall_out_reg_5_NO_SHIFT_REG),
	.data_in(local_bb3_or53_i49),
	.data_out(rnode_1to5_bb3_or53_i49_0_reg_5_NO_SHIFT_REG)
);

defparam rnode_1to5_bb3_or53_i49_0_reg_5_fifo.DEPTH = 5;
defparam rnode_1to5_bb3_or53_i49_0_reg_5_fifo.DATA_WIDTH = 32;
defparam rnode_1to5_bb3_or53_i49_0_reg_5_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_1to5_bb3_or53_i49_0_reg_5_fifo.IMPL = "ll_reg";

assign rnode_1to5_bb3_or53_i49_0_reg_5_inputs_ready_NO_SHIFT_REG = local_bb3_or53_i49_valid_out;
assign local_bb3_or53_i49_stall_in = rnode_1to5_bb3_or53_i49_0_stall_out_reg_5_NO_SHIFT_REG;
assign rnode_1to5_bb3_or53_i49_0_NO_SHIFT_REG = rnode_1to5_bb3_or53_i49_0_reg_5_NO_SHIFT_REG;
assign rnode_1to5_bb3_or53_i49_0_stall_in_reg_5_NO_SHIFT_REG = rnode_1to5_bb3_or53_i49_0_stall_in_NO_SHIFT_REG;
assign rnode_1to5_bb3_or53_i49_0_valid_out_NO_SHIFT_REG = rnode_1to5_bb3_or53_i49_0_valid_out_reg_5_NO_SHIFT_REG;

// Register node:
//  * latency = 1
//  * capacity = 1
 logic rnode_142to143_bb3_or53_i_0_valid_out_NO_SHIFT_REG;
 logic rnode_142to143_bb3_or53_i_0_stall_in_NO_SHIFT_REG;
 logic [31:0] rnode_142to143_bb3_or53_i_0_NO_SHIFT_REG;
 logic rnode_142to143_bb3_or53_i_0_reg_143_inputs_ready_NO_SHIFT_REG;
 logic [31:0] rnode_142to143_bb3_or53_i_0_reg_143_NO_SHIFT_REG;
 logic rnode_142to143_bb3_or53_i_0_valid_out_reg_143_NO_SHIFT_REG;
 logic rnode_142to143_bb3_or53_i_0_stall_in_reg_143_NO_SHIFT_REG;
 logic rnode_142to143_bb3_or53_i_0_stall_out_reg_143_NO_SHIFT_REG;

acl_data_fifo rnode_142to143_bb3_or53_i_0_reg_143_fifo (
	.clock(clock),
	.resetn(resetn),
	.valid_in(rnode_142to143_bb3_or53_i_0_reg_143_inputs_ready_NO_SHIFT_REG),
	.stall_in(rnode_142to143_bb3_or53_i_0_stall_in_reg_143_NO_SHIFT_REG),
	.valid_out(rnode_142to143_bb3_or53_i_0_valid_out_reg_143_NO_SHIFT_REG),
	.stall_out(rnode_142to143_bb3_or53_i_0_stall_out_reg_143_NO_SHIFT_REG),
	.data_in(rnode_1to142_bb3_or53_i_0_NO_SHIFT_REG),
	.data_out(rnode_142to143_bb3_or53_i_0_reg_143_NO_SHIFT_REG)
);

defparam rnode_142to143_bb3_or53_i_0_reg_143_fifo.DEPTH = 2;
defparam rnode_142to143_bb3_or53_i_0_reg_143_fifo.DATA_WIDTH = 32;
defparam rnode_142to143_bb3_or53_i_0_reg_143_fifo.ALLOW_FULL_WRITE = 0;
defparam rnode_142to143_bb3_or53_i_0_reg_143_fifo.IMPL = "ll_reg";

assign rnode_142to143_bb3_or53_i_0_reg_143_inputs_ready_NO_SHIFT_REG = rnode_1to142_bb3_or53_i_0_valid_out_NO_SHIFT_REG;
assign rnode_1to142_bb3_or53_i_0_stall_in_NO_SHIFT_REG = rnode_142to143_bb3_or53_i_0_stall_out_reg_143_NO_SHIFT_REG;
assign rnode_142to143_bb3_or53_i_0_NO_SHIFT_REG = rnode_142to143_bb3_or53_i_0_reg_143_NO_SHIFT_REG;
assign rnode_142to143_bb3_or53_i_0_stall_in_reg_143_NO_SHIFT_REG = rnode_142to143_bb3_or53_i_0_stall_in_NO_SHIFT_REG;
assign rnode_142to143_bb3_or53_i_0_valid_out_NO_SHIFT_REG = rnode_142to143_bb3_or53_i_0_valid_out_reg_143_NO_SHIFT_REG;

// This section implements an unregistered operation.
// 
wire local_bb3_negate_sign14_stall_local;
wire [31:0] local_bb3_negate_sign14;

assign local_bb3_negate_sign14 = (rnode_1to5_bb3_or53_i49_0_NO_SHIFT_REG ^ 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_negate_sign20_stall_local;
wire [31:0] local_bb3_negate_sign20;

assign local_bb3_negate_sign20 = (rnode_142to143_bb3_or53_i_0_NO_SHIFT_REG ^ 32'h80000000);

// This section implements an unregistered operation.
// 
wire local_bb3_cast_after_negation15_stall_local;
wire [31:0] local_bb3_cast_after_negation15;

assign local_bb3_cast_after_negation15 = local_bb3_negate_sign14;

// This section implements an unregistered operation.
// 
wire local_bb3_cast_after_negation21_stall_local;
wire [31:0] local_bb3_cast_after_negation21;

assign local_bb3_cast_after_negation21 = local_bb3_negate_sign20;

// This section implements an unregistered operation.
// 
wire local_bb3_select40_valid_out;
wire local_bb3_select40_stall_in;
wire local_bb3_select40_inputs_ready;
wire local_bb3_select40_stall_local;
wire [31:0] local_bb3_select40;

assign local_bb3_select40_inputs_ready = rnode_1to5_bb3_or53_i49_0_valid_out_NO_SHIFT_REG;
assign local_bb3_select40 = (input_wii_cmp3 ? local_bb3_cast_after_negation15 : 32'h80000000);
assign local_bb3_select40_valid_out = local_bb3_select40_inputs_ready;
assign local_bb3_select40_stall_local = local_bb3_select40_stall_in;
assign rnode_1to5_bb3_or53_i49_0_stall_in_NO_SHIFT_REG = (|local_bb3_select40_stall_local);

// This section implements an unregistered operation.
// 
wire local_bb3_select37_valid_out;
wire local_bb3_select37_stall_in;
wire local_bb3_select37_inputs_ready;
wire local_bb3_select37_stall_local;
wire [31:0] local_bb3_select37;

assign local_bb3_select37_inputs_ready = rnode_142to143_bb3_or53_i_0_valid_out_NO_SHIFT_REG;
assign local_bb3_select37 = (input_wii_cmp3 ? local_bb3_cast_after_negation21 : 32'h80000000);
assign local_bb3_select37_valid_out = local_bb3_select37_inputs_ready;
assign local_bb3_select37_stall_local = local_bb3_select37_stall_in;
assign rnode_142to143_bb3_or53_i_0_stall_in_NO_SHIFT_REG = (|local_bb3_select37_stall_local);

// This section implements a registered operation.
// 
wire local_bb3_st_select40_inputs_ready;
 reg local_bb3_st_select40_valid_out_NO_SHIFT_REG;
wire local_bb3_st_select40_stall_in;
wire local_bb3_st_select40_output_regs_ready;
wire local_bb3_st_select40_fu_stall_out;
wire local_bb3_st_select40_fu_valid_out;
wire [31:0] local_bb3_st_select40_lsu_wackout;
 reg local_bb3_st_select40_NO_SHIFT_REG;
wire local_bb3_st_select40_causedstall;

lsu_top lsu_local_bb3_st_select40 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb3_st_select40_fu_stall_out),
	.i_valid(local_bb3_st_select40_inputs_ready),
	.i_address(rstag_5to5_bb3_arrayidx43),
	.i_writedata(local_bb3_select40),
	.i_cmpdata(),
	.i_predicate(1'b0),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb3_st_select40_output_regs_ready)),
	.o_valid(local_bb3_st_select40_fu_valid_out),
	.o_readdata(),
	.o_input_fifo_depth(),
	.o_writeack(local_bb3_st_select40_lsu_wackout),
	.i_atomic_op(3'h0),
	.o_active(local_bb3_st_select40_active),
	.avm_address(avm_local_bb3_st_select40_address),
	.avm_read(avm_local_bb3_st_select40_read),
	.avm_readdata(avm_local_bb3_st_select40_readdata),
	.avm_write(avm_local_bb3_st_select40_write),
	.avm_writeack(avm_local_bb3_st_select40_writeack),
	.avm_burstcount(avm_local_bb3_st_select40_burstcount),
	.avm_writedata(avm_local_bb3_st_select40_writedata),
	.avm_byteenable(avm_local_bb3_st_select40_byteenable),
	.avm_waitrequest(avm_local_bb3_st_select40_waitrequest),
	.avm_readdatavalid(avm_local_bb3_st_select40_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb3_st_select40.AWIDTH = 30;
defparam lsu_local_bb3_st_select40.WIDTH_BYTES = 4;
defparam lsu_local_bb3_st_select40.MWIDTH_BYTES = 32;
defparam lsu_local_bb3_st_select40.WRITEDATAWIDTH_BYTES = 32;
defparam lsu_local_bb3_st_select40.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb3_st_select40.READ = 0;
defparam lsu_local_bb3_st_select40.ATOMIC = 0;
defparam lsu_local_bb3_st_select40.WIDTH = 32;
defparam lsu_local_bb3_st_select40.MWIDTH = 256;
defparam lsu_local_bb3_st_select40.ATOMIC_WIDTH = 3;
defparam lsu_local_bb3_st_select40.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb3_st_select40.KERNEL_SIDE_MEM_LATENCY = 138;
defparam lsu_local_bb3_st_select40.MEMORY_SIDE_MEM_LATENCY = 10;
defparam lsu_local_bb3_st_select40.USE_WRITE_ACK = 1;
defparam lsu_local_bb3_st_select40.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb3_st_select40.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb3_st_select40.NUMBER_BANKS = 1;
defparam lsu_local_bb3_st_select40.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb3_st_select40.USEINPUTFIFO = 0;
defparam lsu_local_bb3_st_select40.USECACHING = 0;
defparam lsu_local_bb3_st_select40.USEOUTPUTFIFO = 1;
defparam lsu_local_bb3_st_select40.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb3_st_select40.HIGH_FMAX = 1;
defparam lsu_local_bb3_st_select40.ADDRSPACE = 1;
defparam lsu_local_bb3_st_select40.STYLE = "BURST-COALESCED";
defparam lsu_local_bb3_st_select40.USE_BYTE_EN = 0;

assign local_bb3_st_select40_inputs_ready = (local_bb3_select40_valid_out & rstag_5to5_bb3_arrayidx43_valid_out);
assign local_bb3_st_select40_output_regs_ready = (&(~(local_bb3_st_select40_valid_out_NO_SHIFT_REG) | ~(local_bb3_st_select40_stall_in)));
assign local_bb3_select40_stall_in = (local_bb3_st_select40_fu_stall_out | ~(local_bb3_st_select40_inputs_ready));
assign rstag_5to5_bb3_arrayidx43_stall_in = (local_bb3_st_select40_fu_stall_out | ~(local_bb3_st_select40_inputs_ready));
assign local_bb3_st_select40_causedstall = (local_bb3_st_select40_inputs_ready && (local_bb3_st_select40_fu_stall_out && !(~(local_bb3_st_select40_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_st_select40_NO_SHIFT_REG <= 'x;
		local_bb3_st_select40_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_st_select40_output_regs_ready)
		begin
			local_bb3_st_select40_NO_SHIFT_REG <= local_bb3_st_select40_lsu_wackout;
			local_bb3_st_select40_valid_out_NO_SHIFT_REG <= local_bb3_st_select40_fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_st_select40_stall_in))
			begin
				local_bb3_st_select40_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_143to143_bb3_st_select40_valid_out;
wire rstag_143to143_bb3_st_select40_stall_in;
wire rstag_143to143_bb3_st_select40_inputs_ready;
wire rstag_143to143_bb3_st_select40_stall_local;
 reg rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG;
wire rstag_143to143_bb3_st_select40_combined_valid;
 reg rstag_143to143_bb3_st_select40_staging_reg_NO_SHIFT_REG;
wire rstag_143to143_bb3_st_select40;

assign rstag_143to143_bb3_st_select40_inputs_ready = local_bb3_st_select40_valid_out_NO_SHIFT_REG;
assign rstag_143to143_bb3_st_select40 = (rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG ? rstag_143to143_bb3_st_select40_staging_reg_NO_SHIFT_REG : local_bb3_st_select40_NO_SHIFT_REG);
assign rstag_143to143_bb3_st_select40_combined_valid = (rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG | rstag_143to143_bb3_st_select40_inputs_ready);
assign rstag_143to143_bb3_st_select40_valid_out = rstag_143to143_bb3_st_select40_combined_valid;
assign rstag_143to143_bb3_st_select40_stall_local = rstag_143to143_bb3_st_select40_stall_in;
assign local_bb3_st_select40_stall_in = (|rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG <= 1'b0;
		rstag_143to143_bb3_st_select40_staging_reg_NO_SHIFT_REG <= 'x;
	end
	else
	begin
		if (rstag_143to143_bb3_st_select40_stall_local)
		begin
			if (~(rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG))
			begin
				rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG <= rstag_143to143_bb3_st_select40_inputs_ready;
			end
		end
		else
		begin
			rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
		if (~(rstag_143to143_bb3_st_select40_staging_valid_NO_SHIFT_REG))
		begin
			rstag_143to143_bb3_st_select40_staging_reg_NO_SHIFT_REG <= local_bb3_st_select40_NO_SHIFT_REG;
		end
	end
end


// This section implements a registered operation.
// 
wire local_bb3_st_select37_inputs_ready;
 reg local_bb3_st_select37_valid_out_NO_SHIFT_REG;
wire local_bb3_st_select37_stall_in;
wire local_bb3_st_select37_output_regs_ready;
wire local_bb3_st_select37_fu_stall_out;
wire local_bb3_st_select37_fu_valid_out;
wire local_bb3_st_select37_causedstall;

lsu_top lsu_local_bb3_st_select37 (
	.clock(clock),
	.clock2x(clock2x),
	.resetn(resetn),
	.flush(start),
	.stream_base_addr(),
	.stream_size(),
	.stream_reset(),
	.o_stall(local_bb3_st_select37_fu_stall_out),
	.i_valid(local_bb3_st_select37_inputs_ready),
	.i_address(rnode_142to143_bb3_arrayidx48_0_NO_SHIFT_REG),
	.i_writedata(local_bb3_select37),
	.i_cmpdata(),
	.i_predicate(1'b0),
	.i_bitwiseor(64'h0),
	.i_byteenable(),
	.i_stall(~(local_bb3_st_select37_output_regs_ready)),
	.o_valid(local_bb3_st_select37_fu_valid_out),
	.o_readdata(),
	.o_input_fifo_depth(),
	.o_writeack(),
	.i_atomic_op(3'h0),
	.o_active(local_bb3_st_select37_active),
	.avm_address(avm_local_bb3_st_select37_address),
	.avm_read(avm_local_bb3_st_select37_read),
	.avm_readdata(avm_local_bb3_st_select37_readdata),
	.avm_write(avm_local_bb3_st_select37_write),
	.avm_writeack(avm_local_bb3_st_select37_writeack),
	.avm_burstcount(avm_local_bb3_st_select37_burstcount),
	.avm_writedata(avm_local_bb3_st_select37_writedata),
	.avm_byteenable(avm_local_bb3_st_select37_byteenable),
	.avm_waitrequest(avm_local_bb3_st_select37_waitrequest),
	.avm_readdatavalid(avm_local_bb3_st_select37_readdatavalid),
	.profile_bw(),
	.profile_bw_incr(),
	.profile_total_ivalid(),
	.profile_total_req(),
	.profile_i_stall_count(),
	.profile_o_stall_count(),
	.profile_avm_readwrite_count(),
	.profile_avm_burstcount_total(),
	.profile_avm_burstcount_total_incr(),
	.profile_req_cache_hit_count(),
	.profile_extra_unaligned_reqs(),
	.profile_avm_stall()
);

defparam lsu_local_bb3_st_select37.AWIDTH = 30;
defparam lsu_local_bb3_st_select37.WIDTH_BYTES = 4;
defparam lsu_local_bb3_st_select37.MWIDTH_BYTES = 32;
defparam lsu_local_bb3_st_select37.WRITEDATAWIDTH_BYTES = 32;
defparam lsu_local_bb3_st_select37.ALIGNMENT_BYTES = 4;
defparam lsu_local_bb3_st_select37.READ = 0;
defparam lsu_local_bb3_st_select37.ATOMIC = 0;
defparam lsu_local_bb3_st_select37.WIDTH = 32;
defparam lsu_local_bb3_st_select37.MWIDTH = 256;
defparam lsu_local_bb3_st_select37.ATOMIC_WIDTH = 3;
defparam lsu_local_bb3_st_select37.BURSTCOUNT_WIDTH = 5;
defparam lsu_local_bb3_st_select37.KERNEL_SIDE_MEM_LATENCY = 4;
defparam lsu_local_bb3_st_select37.MEMORY_SIDE_MEM_LATENCY = 10;
defparam lsu_local_bb3_st_select37.USE_WRITE_ACK = 0;
defparam lsu_local_bb3_st_select37.ENABLE_BANKED_MEMORY = 0;
defparam lsu_local_bb3_st_select37.ABITS_PER_LMEM_BANK = 0;
defparam lsu_local_bb3_st_select37.NUMBER_BANKS = 1;
defparam lsu_local_bb3_st_select37.LMEM_ADDR_PERMUTATION_STYLE = 0;
defparam lsu_local_bb3_st_select37.USEINPUTFIFO = 0;
defparam lsu_local_bb3_st_select37.USECACHING = 0;
defparam lsu_local_bb3_st_select37.USEOUTPUTFIFO = 1;
defparam lsu_local_bb3_st_select37.FORCE_NOP_SUPPORT = 0;
defparam lsu_local_bb3_st_select37.HIGH_FMAX = 1;
defparam lsu_local_bb3_st_select37.ADDRSPACE = 1;
defparam lsu_local_bb3_st_select37.STYLE = "BURST-COALESCED";
defparam lsu_local_bb3_st_select37.USE_BYTE_EN = 0;

assign local_bb3_st_select37_inputs_ready = (local_bb3_select37_valid_out & rnode_142to143_bb3_arrayidx48_0_valid_out_NO_SHIFT_REG & rstag_143to143_bb3_st_select40_valid_out);
assign local_bb3_st_select37_output_regs_ready = (&(~(local_bb3_st_select37_valid_out_NO_SHIFT_REG) | ~(local_bb3_st_select37_stall_in)));
assign local_bb3_select37_stall_in = (local_bb3_st_select37_fu_stall_out | ~(local_bb3_st_select37_inputs_ready));
assign rnode_142to143_bb3_arrayidx48_0_stall_in_NO_SHIFT_REG = (local_bb3_st_select37_fu_stall_out | ~(local_bb3_st_select37_inputs_ready));
assign rstag_143to143_bb3_st_select40_stall_in = (local_bb3_st_select37_fu_stall_out | ~(local_bb3_st_select37_inputs_ready));
assign local_bb3_st_select37_causedstall = (local_bb3_st_select37_inputs_ready && (local_bb3_st_select37_fu_stall_out && !(~(local_bb3_st_select37_output_regs_ready))));

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		local_bb3_st_select37_valid_out_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (local_bb3_st_select37_output_regs_ready)
		begin
			local_bb3_st_select37_valid_out_NO_SHIFT_REG <= local_bb3_st_select37_fu_valid_out;
		end
		else
		begin
			if (~(local_bb3_st_select37_stall_in))
			begin
				local_bb3_st_select37_valid_out_NO_SHIFT_REG <= 1'b0;
			end
		end
	end
end


// This section implements a staging register.
// 
wire rstag_147to147_bb3_st_select37_valid_out;
wire rstag_147to147_bb3_st_select37_stall_in;
wire rstag_147to147_bb3_st_select37_inputs_ready;
wire rstag_147to147_bb3_st_select37_stall_local;
 reg rstag_147to147_bb3_st_select37_staging_valid_NO_SHIFT_REG;
wire rstag_147to147_bb3_st_select37_combined_valid;

assign rstag_147to147_bb3_st_select37_inputs_ready = local_bb3_st_select37_valid_out_NO_SHIFT_REG;
assign rstag_147to147_bb3_st_select37_combined_valid = (rstag_147to147_bb3_st_select37_staging_valid_NO_SHIFT_REG | rstag_147to147_bb3_st_select37_inputs_ready);
assign rstag_147to147_bb3_st_select37_valid_out = rstag_147to147_bb3_st_select37_combined_valid;
assign rstag_147to147_bb3_st_select37_stall_local = rstag_147to147_bb3_st_select37_stall_in;
assign local_bb3_st_select37_stall_in = (|rstag_147to147_bb3_st_select37_staging_valid_NO_SHIFT_REG);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		rstag_147to147_bb3_st_select37_staging_valid_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		if (rstag_147to147_bb3_st_select37_stall_local)
		begin
			if (~(rstag_147to147_bb3_st_select37_staging_valid_NO_SHIFT_REG))
			begin
				rstag_147to147_bb3_st_select37_staging_valid_NO_SHIFT_REG <= rstag_147to147_bb3_st_select37_inputs_ready;
			end
		end
		else
		begin
			rstag_147to147_bb3_st_select37_staging_valid_NO_SHIFT_REG <= 1'b0;
		end
	end
end


// This section describes the behaviour of the BRANCH node.
wire branch_var__inputs_ready;
wire branch_var__output_regs_ready;

assign branch_var__inputs_ready = rstag_147to147_bb3_st_select37_valid_out;
assign branch_var__output_regs_ready = ~(stall_in);
assign rstag_147to147_bb3_st_select37_stall_in = (~(branch_var__output_regs_ready) | ~(branch_var__inputs_ready));
assign valid_out = branch_var__inputs_ready;

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

module Matmul_function
	(
		input 		clock,
		input 		resetn,
		input [31:0] 		input_global_id_0,
		input [31:0] 		input_global_id_1,
		output 		stall_out,
		input 		valid_in,
		output 		valid_out,
		input 		stall_in,
		input [31:0] 		workgroup_size,
		input [255:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_readdata,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_readdatavalid,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_waitrequest,
		output [29:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_address,
		output 		avm_local_bb2_ld_memcoalesce_m1r_load_0_read,
		output 		avm_local_bb2_ld_memcoalesce_m1r_load_0_write,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_writeack,
		output [255:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_writedata,
		output [31:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_byteenable,
		output [4:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_burstcount,
		input [255:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_readdata,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_readdatavalid,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_waitrequest,
		output [29:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_address,
		output 		avm_local_bb2_ld_memcoalesce_m1i_load_0_read,
		output 		avm_local_bb2_ld_memcoalesce_m1i_load_0_write,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_writeack,
		output [255:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_writedata,
		output [31:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_byteenable,
		output [4:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_burstcount,
		input [255:0] 		avm_local_bb2_ld__readdata,
		input 		avm_local_bb2_ld__readdatavalid,
		input 		avm_local_bb2_ld__waitrequest,
		output [29:0] 		avm_local_bb2_ld__address,
		output 		avm_local_bb2_ld__read,
		output 		avm_local_bb2_ld__write,
		input 		avm_local_bb2_ld__writeack,
		output [255:0] 		avm_local_bb2_ld__writedata,
		output [31:0] 		avm_local_bb2_ld__byteenable,
		output [4:0] 		avm_local_bb2_ld__burstcount,
		input [255:0] 		avm_local_bb2_ld__u1_readdata,
		input 		avm_local_bb2_ld__u1_readdatavalid,
		input 		avm_local_bb2_ld__u1_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u1_address,
		output 		avm_local_bb2_ld__u1_read,
		output 		avm_local_bb2_ld__u1_write,
		input 		avm_local_bb2_ld__u1_writeack,
		output [255:0] 		avm_local_bb2_ld__u1_writedata,
		output [31:0] 		avm_local_bb2_ld__u1_byteenable,
		output [4:0] 		avm_local_bb2_ld__u1_burstcount,
		input [255:0] 		avm_local_bb2_ld__u2_readdata,
		input 		avm_local_bb2_ld__u2_readdatavalid,
		input 		avm_local_bb2_ld__u2_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u2_address,
		output 		avm_local_bb2_ld__u2_read,
		output 		avm_local_bb2_ld__u2_write,
		input 		avm_local_bb2_ld__u2_writeack,
		output [255:0] 		avm_local_bb2_ld__u2_writedata,
		output [31:0] 		avm_local_bb2_ld__u2_byteenable,
		output [4:0] 		avm_local_bb2_ld__u2_burstcount,
		input [255:0] 		avm_local_bb2_ld__u3_readdata,
		input 		avm_local_bb2_ld__u3_readdatavalid,
		input 		avm_local_bb2_ld__u3_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u3_address,
		output 		avm_local_bb2_ld__u3_read,
		output 		avm_local_bb2_ld__u3_write,
		input 		avm_local_bb2_ld__u3_writeack,
		output [255:0] 		avm_local_bb2_ld__u3_writedata,
		output [31:0] 		avm_local_bb2_ld__u3_byteenable,
		output [4:0] 		avm_local_bb2_ld__u3_burstcount,
		input [255:0] 		avm_local_bb3_st_select40_readdata,
		input 		avm_local_bb3_st_select40_readdatavalid,
		input 		avm_local_bb3_st_select40_waitrequest,
		output [29:0] 		avm_local_bb3_st_select40_address,
		output 		avm_local_bb3_st_select40_read,
		output 		avm_local_bb3_st_select40_write,
		input 		avm_local_bb3_st_select40_writeack,
		output [255:0] 		avm_local_bb3_st_select40_writedata,
		output [31:0] 		avm_local_bb3_st_select40_byteenable,
		output [4:0] 		avm_local_bb3_st_select40_burstcount,
		input [255:0] 		avm_local_bb3_st_select37_readdata,
		input 		avm_local_bb3_st_select37_readdatavalid,
		input 		avm_local_bb3_st_select37_waitrequest,
		output [29:0] 		avm_local_bb3_st_select37_address,
		output 		avm_local_bb3_st_select37_read,
		output 		avm_local_bb3_st_select37_write,
		input 		avm_local_bb3_st_select37_writeack,
		output [255:0] 		avm_local_bb3_st_select37_writedata,
		output [31:0] 		avm_local_bb3_st_select37_byteenable,
		output [4:0] 		avm_local_bb3_st_select37_burstcount,
		input 		start,
		input [31:0] 		input_c1f2,
		input 		clock2x,
		input [63:0] 		input_m1r,
		input [63:0] 		input_m1i,
		input [31:0] 		input_col_m2,
		input [63:0] 		input_m2r,
		input [63:0] 		input_m2i,
		input [63:0] 		input_rer,
		input [63:0] 		input_rei,
		output reg 		has_a_write_pending,
		output reg 		has_a_lsu_active
	);


wire [31:0] cur_cycle;
wire bb_0_stall_out;
wire bb_0_valid_out;
wire bb_0_lvb_bb0_cmp3;
wire bb_0_lvb_bb0_cmp3_NEG;
wire [31:0] bb_0_lvb_input_global_id_0;
wire [31:0] bb_0_lvb_input_global_id_1;
wire bb_1_stall_out;
wire bb_1_valid_out;
wire [63:0] bb_1_lvb_bb1_var_;
wire [31:0] bb_1_lvb_input_global_id_0;
wire [31:0] bb_1_lvb_input_global_id_1;
wire bb_2_stall_out_0;
wire bb_2_stall_out_1;
wire bb_2_valid_out_0;
wire [63:0] bb_2_lvb_var__0;
wire [63:0] bb_2_lvb_bb2_indvars_iv_next_1_0;
wire bb_2_lvb_bb2_exitcond_0;
wire [159:0] bb_2_lvb_bb2_c0_exit_c0_exi4_0;
wire [31:0] bb_2_lvb_bb2_c0_exe3_0;
wire [31:0] bb_2_lvb_bb2_c0_exe4_0;
wire [31:0] bb_2_lvb_input_global_id_0_0;
wire [31:0] bb_2_lvb_input_global_id_1_0;
wire bb_2_valid_out_1;
wire [63:0] bb_2_lvb_var__1;
wire [63:0] bb_2_lvb_bb2_indvars_iv_next_1_1;
wire bb_2_lvb_bb2_exitcond_1;
wire [159:0] bb_2_lvb_bb2_c0_exit_c0_exi4_1;
wire [31:0] bb_2_lvb_bb2_c0_exe3_1;
wire [31:0] bb_2_lvb_bb2_c0_exe4_1;
wire [31:0] bb_2_lvb_input_global_id_0_1;
wire [31:0] bb_2_lvb_input_global_id_1_1;
wire bb_2_local_bb2_ld_memcoalesce_m1r_load_0_active;
wire bb_2_local_bb2_ld_memcoalesce_m1i_load_0_active;
wire bb_2_local_bb2_ld__active;
wire bb_2_local_bb2_ld__u1_active;
wire bb_2_local_bb2_ld__u2_active;
wire bb_2_local_bb2_ld__u3_active;
wire bb_3_stall_out;
wire bb_3_valid_out;
wire bb_3_local_bb3_st_select40_active;
wire bb_3_local_bb3_st_select37_active;
wire loop_limiter_0_stall_out;
wire loop_limiter_0_valid_out;
wire [1:0] writes_pending;
wire [7:0] lsus_active;

Matmul_basic_block_0 Matmul_basic_block_0 (
	.clock(clock),
	.resetn(resetn),
	.start(start),
	.input_c1f2(input_c1f2),
	.valid_in(valid_in),
	.stall_out(bb_0_stall_out),
	.input_global_id_0(input_global_id_0),
	.input_global_id_1(input_global_id_1),
	.valid_out(bb_0_valid_out),
	.stall_in(bb_1_stall_out),
	.lvb_bb0_cmp3(bb_0_lvb_bb0_cmp3),
	.lvb_bb0_cmp3_NEG(bb_0_lvb_bb0_cmp3_NEG),
	.lvb_input_global_id_0(bb_0_lvb_input_global_id_0),
	.lvb_input_global_id_1(bb_0_lvb_input_global_id_1),
	.workgroup_size(workgroup_size)
);


Matmul_basic_block_1 Matmul_basic_block_1 (
	.clock(clock),
	.resetn(resetn),
	.input_c1f2(input_c1f2),
	.input_wii_cmp3(bb_0_lvb_bb0_cmp3),
	.input_wii_cmp3_NEG(bb_0_lvb_bb0_cmp3_NEG),
	.valid_in(bb_0_valid_out),
	.stall_out(bb_1_stall_out),
	.input_global_id_0(bb_0_lvb_input_global_id_0),
	.input_global_id_1(bb_0_lvb_input_global_id_1),
	.valid_out(bb_1_valid_out),
	.stall_in(loop_limiter_0_stall_out),
	.lvb_bb1_var_(bb_1_lvb_bb1_var_),
	.lvb_input_global_id_0(bb_1_lvb_input_global_id_0),
	.lvb_input_global_id_1(bb_1_lvb_input_global_id_1),
	.workgroup_size(workgroup_size),
	.start(start)
);


Matmul_basic_block_2 Matmul_basic_block_2 (
	.clock(clock),
	.resetn(resetn),
	.input_m1r(input_m1r),
	.input_m1i(input_m1i),
	.input_col_m2(input_col_m2),
	.input_c1f2(input_c1f2),
	.input_m2r(input_m2r),
	.input_m2i(input_m2i),
	.input_wii_cmp3(bb_0_lvb_bb0_cmp3),
	.input_wii_cmp3_NEG(bb_0_lvb_bb0_cmp3_NEG),
	.valid_in_0(bb_2_valid_out_1),
	.stall_out_0(bb_2_stall_out_0),
	.input_var__0(bb_2_lvb_var__1),
	.input_indvars_iv_0(bb_2_lvb_bb2_indvars_iv_next_1_1),
	.input_tmpi_06_0(bb_2_lvb_bb2_c0_exe4_1),
	.input_tmpr_05_0(bb_2_lvb_bb2_c0_exe3_1),
	.input_global_id_0_0(bb_2_lvb_input_global_id_0_1),
	.input_global_id_1_0(bb_2_lvb_input_global_id_1_1),
	.valid_in_1(loop_limiter_0_valid_out),
	.stall_out_1(bb_2_stall_out_1),
	.input_var__1(bb_1_lvb_bb1_var_),
	.input_indvars_iv_1(64'h0),
	.input_tmpi_06_1(32'h0),
	.input_tmpr_05_1(32'h0),
	.input_global_id_0_1(bb_1_lvb_input_global_id_0),
	.input_global_id_1_1(bb_1_lvb_input_global_id_1),
	.valid_out_0(bb_2_valid_out_0),
	.stall_in_0(bb_3_stall_out),
	.lvb_var__0(bb_2_lvb_var__0),
	.lvb_bb2_indvars_iv_next_1_0(bb_2_lvb_bb2_indvars_iv_next_1_0),
	.lvb_bb2_exitcond_0(bb_2_lvb_bb2_exitcond_0),
	.lvb_bb2_c0_exit_c0_exi4_0(bb_2_lvb_bb2_c0_exit_c0_exi4_0),
	.lvb_bb2_c0_exe3_0(bb_2_lvb_bb2_c0_exe3_0),
	.lvb_bb2_c0_exe4_0(bb_2_lvb_bb2_c0_exe4_0),
	.lvb_input_global_id_0_0(bb_2_lvb_input_global_id_0_0),
	.lvb_input_global_id_1_0(bb_2_lvb_input_global_id_1_0),
	.valid_out_1(bb_2_valid_out_1),
	.stall_in_1(bb_2_stall_out_0),
	.lvb_var__1(bb_2_lvb_var__1),
	.lvb_bb2_indvars_iv_next_1_1(bb_2_lvb_bb2_indvars_iv_next_1_1),
	.lvb_bb2_exitcond_1(bb_2_lvb_bb2_exitcond_1),
	.lvb_bb2_c0_exit_c0_exi4_1(bb_2_lvb_bb2_c0_exit_c0_exi4_1),
	.lvb_bb2_c0_exe3_1(bb_2_lvb_bb2_c0_exe3_1),
	.lvb_bb2_c0_exe4_1(bb_2_lvb_bb2_c0_exe4_1),
	.lvb_input_global_id_0_1(bb_2_lvb_input_global_id_0_1),
	.lvb_input_global_id_1_1(bb_2_lvb_input_global_id_1_1),
	.workgroup_size(workgroup_size),
	.start(start),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_readdata(avm_local_bb2_ld_memcoalesce_m1r_load_0_readdata),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_readdatavalid(avm_local_bb2_ld_memcoalesce_m1r_load_0_readdatavalid),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_waitrequest(avm_local_bb2_ld_memcoalesce_m1r_load_0_waitrequest),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_address(avm_local_bb2_ld_memcoalesce_m1r_load_0_address),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_read(avm_local_bb2_ld_memcoalesce_m1r_load_0_read),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_write(avm_local_bb2_ld_memcoalesce_m1r_load_0_write),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_writeack(avm_local_bb2_ld_memcoalesce_m1r_load_0_writeack),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_writedata(avm_local_bb2_ld_memcoalesce_m1r_load_0_writedata),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_byteenable(avm_local_bb2_ld_memcoalesce_m1r_load_0_byteenable),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_burstcount(avm_local_bb2_ld_memcoalesce_m1r_load_0_burstcount),
	.local_bb2_ld_memcoalesce_m1r_load_0_active(bb_2_local_bb2_ld_memcoalesce_m1r_load_0_active),
	.clock2x(clock2x),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_readdata(avm_local_bb2_ld_memcoalesce_m1i_load_0_readdata),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_readdatavalid(avm_local_bb2_ld_memcoalesce_m1i_load_0_readdatavalid),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_waitrequest(avm_local_bb2_ld_memcoalesce_m1i_load_0_waitrequest),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_address(avm_local_bb2_ld_memcoalesce_m1i_load_0_address),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_read(avm_local_bb2_ld_memcoalesce_m1i_load_0_read),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_write(avm_local_bb2_ld_memcoalesce_m1i_load_0_write),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_writeack(avm_local_bb2_ld_memcoalesce_m1i_load_0_writeack),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_writedata(avm_local_bb2_ld_memcoalesce_m1i_load_0_writedata),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_byteenable(avm_local_bb2_ld_memcoalesce_m1i_load_0_byteenable),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_burstcount(avm_local_bb2_ld_memcoalesce_m1i_load_0_burstcount),
	.local_bb2_ld_memcoalesce_m1i_load_0_active(bb_2_local_bb2_ld_memcoalesce_m1i_load_0_active),
	.avm_local_bb2_ld__readdata(avm_local_bb2_ld__readdata),
	.avm_local_bb2_ld__readdatavalid(avm_local_bb2_ld__readdatavalid),
	.avm_local_bb2_ld__waitrequest(avm_local_bb2_ld__waitrequest),
	.avm_local_bb2_ld__address(avm_local_bb2_ld__address),
	.avm_local_bb2_ld__read(avm_local_bb2_ld__read),
	.avm_local_bb2_ld__write(avm_local_bb2_ld__write),
	.avm_local_bb2_ld__writeack(avm_local_bb2_ld__writeack),
	.avm_local_bb2_ld__writedata(avm_local_bb2_ld__writedata),
	.avm_local_bb2_ld__byteenable(avm_local_bb2_ld__byteenable),
	.avm_local_bb2_ld__burstcount(avm_local_bb2_ld__burstcount),
	.local_bb2_ld__active(bb_2_local_bb2_ld__active),
	.avm_local_bb2_ld__u1_readdata(avm_local_bb2_ld__u1_readdata),
	.avm_local_bb2_ld__u1_readdatavalid(avm_local_bb2_ld__u1_readdatavalid),
	.avm_local_bb2_ld__u1_waitrequest(avm_local_bb2_ld__u1_waitrequest),
	.avm_local_bb2_ld__u1_address(avm_local_bb2_ld__u1_address),
	.avm_local_bb2_ld__u1_read(avm_local_bb2_ld__u1_read),
	.avm_local_bb2_ld__u1_write(avm_local_bb2_ld__u1_write),
	.avm_local_bb2_ld__u1_writeack(avm_local_bb2_ld__u1_writeack),
	.avm_local_bb2_ld__u1_writedata(avm_local_bb2_ld__u1_writedata),
	.avm_local_bb2_ld__u1_byteenable(avm_local_bb2_ld__u1_byteenable),
	.avm_local_bb2_ld__u1_burstcount(avm_local_bb2_ld__u1_burstcount),
	.local_bb2_ld__u1_active(bb_2_local_bb2_ld__u1_active),
	.avm_local_bb2_ld__u2_readdata(avm_local_bb2_ld__u2_readdata),
	.avm_local_bb2_ld__u2_readdatavalid(avm_local_bb2_ld__u2_readdatavalid),
	.avm_local_bb2_ld__u2_waitrequest(avm_local_bb2_ld__u2_waitrequest),
	.avm_local_bb2_ld__u2_address(avm_local_bb2_ld__u2_address),
	.avm_local_bb2_ld__u2_read(avm_local_bb2_ld__u2_read),
	.avm_local_bb2_ld__u2_write(avm_local_bb2_ld__u2_write),
	.avm_local_bb2_ld__u2_writeack(avm_local_bb2_ld__u2_writeack),
	.avm_local_bb2_ld__u2_writedata(avm_local_bb2_ld__u2_writedata),
	.avm_local_bb2_ld__u2_byteenable(avm_local_bb2_ld__u2_byteenable),
	.avm_local_bb2_ld__u2_burstcount(avm_local_bb2_ld__u2_burstcount),
	.local_bb2_ld__u2_active(bb_2_local_bb2_ld__u2_active),
	.avm_local_bb2_ld__u3_readdata(avm_local_bb2_ld__u3_readdata),
	.avm_local_bb2_ld__u3_readdatavalid(avm_local_bb2_ld__u3_readdatavalid),
	.avm_local_bb2_ld__u3_waitrequest(avm_local_bb2_ld__u3_waitrequest),
	.avm_local_bb2_ld__u3_address(avm_local_bb2_ld__u3_address),
	.avm_local_bb2_ld__u3_read(avm_local_bb2_ld__u3_read),
	.avm_local_bb2_ld__u3_write(avm_local_bb2_ld__u3_write),
	.avm_local_bb2_ld__u3_writeack(avm_local_bb2_ld__u3_writeack),
	.avm_local_bb2_ld__u3_writedata(avm_local_bb2_ld__u3_writedata),
	.avm_local_bb2_ld__u3_byteenable(avm_local_bb2_ld__u3_byteenable),
	.avm_local_bb2_ld__u3_burstcount(avm_local_bb2_ld__u3_burstcount),
	.local_bb2_ld__u3_active(bb_2_local_bb2_ld__u3_active)
);


Matmul_basic_block_3 Matmul_basic_block_3 (
	.clock(clock),
	.resetn(resetn),
	.input_col_m2(input_col_m2),
	.input_rer(input_rer),
	.input_rei(input_rei),
	.input_wii_cmp3(bb_0_lvb_bb0_cmp3),
	.valid_in(bb_2_valid_out_0),
	.stall_out(bb_3_stall_out),
	.input_exitcond(bb_2_lvb_bb2_exitcond_0),
	.input_c0_exit_c0_exi4(bb_2_lvb_bb2_c0_exit_c0_exi4_0),
	.input_c0_exe3(bb_2_lvb_bb2_c0_exe3_0),
	.input_c0_exe4(bb_2_lvb_bb2_c0_exe4_0),
	.input_global_id_0(bb_2_lvb_input_global_id_0_0),
	.input_global_id_1(bb_2_lvb_input_global_id_1_0),
	.valid_out(bb_3_valid_out),
	.stall_in(stall_in),
	.workgroup_size(workgroup_size),
	.start(start),
	.avm_local_bb3_st_select40_readdata(avm_local_bb3_st_select40_readdata),
	.avm_local_bb3_st_select40_readdatavalid(avm_local_bb3_st_select40_readdatavalid),
	.avm_local_bb3_st_select40_waitrequest(avm_local_bb3_st_select40_waitrequest),
	.avm_local_bb3_st_select40_address(avm_local_bb3_st_select40_address),
	.avm_local_bb3_st_select40_read(avm_local_bb3_st_select40_read),
	.avm_local_bb3_st_select40_write(avm_local_bb3_st_select40_write),
	.avm_local_bb3_st_select40_writeack(avm_local_bb3_st_select40_writeack),
	.avm_local_bb3_st_select40_writedata(avm_local_bb3_st_select40_writedata),
	.avm_local_bb3_st_select40_byteenable(avm_local_bb3_st_select40_byteenable),
	.avm_local_bb3_st_select40_burstcount(avm_local_bb3_st_select40_burstcount),
	.local_bb3_st_select40_active(bb_3_local_bb3_st_select40_active),
	.clock2x(clock2x),
	.avm_local_bb3_st_select37_readdata(avm_local_bb3_st_select37_readdata),
	.avm_local_bb3_st_select37_readdatavalid(avm_local_bb3_st_select37_readdatavalid),
	.avm_local_bb3_st_select37_waitrequest(avm_local_bb3_st_select37_waitrequest),
	.avm_local_bb3_st_select37_address(avm_local_bb3_st_select37_address),
	.avm_local_bb3_st_select37_read(avm_local_bb3_st_select37_read),
	.avm_local_bb3_st_select37_write(avm_local_bb3_st_select37_write),
	.avm_local_bb3_st_select37_writeack(avm_local_bb3_st_select37_writeack),
	.avm_local_bb3_st_select37_writedata(avm_local_bb3_st_select37_writedata),
	.avm_local_bb3_st_select37_byteenable(avm_local_bb3_st_select37_byteenable),
	.avm_local_bb3_st_select37_burstcount(avm_local_bb3_st_select37_burstcount),
	.local_bb3_st_select37_active(bb_3_local_bb3_st_select37_active)
);


acl_loop_limiter loop_limiter_0 (
	.clock(clock),
	.resetn(resetn),
	.i_valid(bb_1_valid_out),
	.i_stall(bb_2_stall_out_1),
	.i_valid_exit(bb_2_valid_out_0),
	.i_stall_exit(bb_3_stall_out),
	.o_valid(loop_limiter_0_valid_out),
	.o_stall(loop_limiter_0_stall_out)
);

defparam loop_limiter_0.ENTRY_WIDTH = 1;
defparam loop_limiter_0.EXIT_WIDTH = 1;
defparam loop_limiter_0.THRESHOLD = 197;

Matmul_sys_cycle_time system_cycle_time_module (
	.clock(clock),
	.resetn(resetn),
	.cur_cycle(cur_cycle)
);


assign valid_out = bb_3_valid_out;
assign stall_out = bb_0_stall_out;
assign writes_pending[0] = bb_3_local_bb3_st_select40_active;
assign writes_pending[1] = bb_3_local_bb3_st_select37_active;
assign lsus_active[0] = bb_2_local_bb2_ld_memcoalesce_m1r_load_0_active;
assign lsus_active[1] = bb_2_local_bb2_ld_memcoalesce_m1i_load_0_active;
assign lsus_active[2] = bb_2_local_bb2_ld__active;
assign lsus_active[3] = bb_2_local_bb2_ld__u1_active;
assign lsus_active[4] = bb_2_local_bb2_ld__u2_active;
assign lsus_active[5] = bb_2_local_bb2_ld__u3_active;
assign lsus_active[6] = bb_3_local_bb3_st_select40_active;
assign lsus_active[7] = bb_3_local_bb3_st_select37_active;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		has_a_write_pending <= 1'b0;
		has_a_lsu_active <= 1'b0;
	end
	else
	begin
		has_a_write_pending <= (|writes_pending);
		has_a_lsu_active <= (|lsus_active);
	end
end

endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

module Matmul_function_wrapper
	(
		input 		clock,
		input 		resetn,
		input 		clock2x,
		input 		local_router_hang,
		input 		avs_cra_read,
		input 		avs_cra_write,
		input [4:0] 		avs_cra_address,
		input [63:0] 		avs_cra_writedata,
		input [7:0] 		avs_cra_byteenable,
		output 		avs_cra_waitrequest,
		output reg [63:0] 		avs_cra_readdata,
		output reg 		avs_cra_readdatavalid,
		output 		cra_irq,
		input [255:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_readdata,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_readdatavalid,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_waitrequest,
		output [29:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_address,
		output 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_read,
		output 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_write,
		input 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_writeack,
		output [255:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_writedata,
		output [31:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_burstcount,
		input [255:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_readdata,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_readdatavalid,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_waitrequest,
		output [29:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_address,
		output 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_read,
		output 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_write,
		input 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_writeack,
		output [255:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_writedata,
		output [31:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_burstcount,
		input [255:0] 		avm_local_bb2_ld__inst0_readdata,
		input 		avm_local_bb2_ld__inst0_readdatavalid,
		input 		avm_local_bb2_ld__inst0_waitrequest,
		output [29:0] 		avm_local_bb2_ld__inst0_address,
		output 		avm_local_bb2_ld__inst0_read,
		output 		avm_local_bb2_ld__inst0_write,
		input 		avm_local_bb2_ld__inst0_writeack,
		output [255:0] 		avm_local_bb2_ld__inst0_writedata,
		output [31:0] 		avm_local_bb2_ld__inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld__inst0_burstcount,
		input [255:0] 		avm_local_bb2_ld__u1_inst0_readdata,
		input 		avm_local_bb2_ld__u1_inst0_readdatavalid,
		input 		avm_local_bb2_ld__u1_inst0_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u1_inst0_address,
		output 		avm_local_bb2_ld__u1_inst0_read,
		output 		avm_local_bb2_ld__u1_inst0_write,
		input 		avm_local_bb2_ld__u1_inst0_writeack,
		output [255:0] 		avm_local_bb2_ld__u1_inst0_writedata,
		output [31:0] 		avm_local_bb2_ld__u1_inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld__u1_inst0_burstcount,
		input [255:0] 		avm_local_bb2_ld__u2_inst0_readdata,
		input 		avm_local_bb2_ld__u2_inst0_readdatavalid,
		input 		avm_local_bb2_ld__u2_inst0_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u2_inst0_address,
		output 		avm_local_bb2_ld__u2_inst0_read,
		output 		avm_local_bb2_ld__u2_inst0_write,
		input 		avm_local_bb2_ld__u2_inst0_writeack,
		output [255:0] 		avm_local_bb2_ld__u2_inst0_writedata,
		output [31:0] 		avm_local_bb2_ld__u2_inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld__u2_inst0_burstcount,
		input [255:0] 		avm_local_bb2_ld__u3_inst0_readdata,
		input 		avm_local_bb2_ld__u3_inst0_readdatavalid,
		input 		avm_local_bb2_ld__u3_inst0_waitrequest,
		output [29:0] 		avm_local_bb2_ld__u3_inst0_address,
		output 		avm_local_bb2_ld__u3_inst0_read,
		output 		avm_local_bb2_ld__u3_inst0_write,
		input 		avm_local_bb2_ld__u3_inst0_writeack,
		output [255:0] 		avm_local_bb2_ld__u3_inst0_writedata,
		output [31:0] 		avm_local_bb2_ld__u3_inst0_byteenable,
		output [4:0] 		avm_local_bb2_ld__u3_inst0_burstcount,
		input [255:0] 		avm_local_bb3_st_select40_inst0_readdata,
		input 		avm_local_bb3_st_select40_inst0_readdatavalid,
		input 		avm_local_bb3_st_select40_inst0_waitrequest,
		output [29:0] 		avm_local_bb3_st_select40_inst0_address,
		output 		avm_local_bb3_st_select40_inst0_read,
		output 		avm_local_bb3_st_select40_inst0_write,
		input 		avm_local_bb3_st_select40_inst0_writeack,
		output [255:0] 		avm_local_bb3_st_select40_inst0_writedata,
		output [31:0] 		avm_local_bb3_st_select40_inst0_byteenable,
		output [4:0] 		avm_local_bb3_st_select40_inst0_burstcount,
		input [255:0] 		avm_local_bb3_st_select37_inst0_readdata,
		input 		avm_local_bb3_st_select37_inst0_readdatavalid,
		input 		avm_local_bb3_st_select37_inst0_waitrequest,
		output [29:0] 		avm_local_bb3_st_select37_inst0_address,
		output 		avm_local_bb3_st_select37_inst0_read,
		output 		avm_local_bb3_st_select37_inst0_write,
		input 		avm_local_bb3_st_select37_inst0_writeack,
		output [255:0] 		avm_local_bb3_st_select37_inst0_writedata,
		output [31:0] 		avm_local_bb3_st_select37_inst0_byteenable,
		output [4:0] 		avm_local_bb3_st_select37_inst0_burstcount
	);

// Responsible for interfacing a kernel with the outside world. It comprises a
// slave interface to specify the kernel arguments and retain kernel status. 

// This section of the wrapper implements the slave interface.
// twoXclock_consumer uses clock2x, even if nobody inside the kernel does. Keeps interface to acl_iface consistent for all kernels.
 reg start_NO_SHIFT_REG;
 reg started_NO_SHIFT_REG;
wire finish;
 reg [31:0] status_NO_SHIFT_REG;
wire has_a_write_pending;
wire has_a_lsu_active;
 reg [447:0] kernel_arguments_NO_SHIFT_REG;
 reg twoXclock_consumer_NO_SHIFT_REG /* synthesis  preserve  noprune  */;
 reg [31:0] workgroup_size_NO_SHIFT_REG;
 reg [31:0] global_size_NO_SHIFT_REG[2:0];
 reg [31:0] num_groups_NO_SHIFT_REG[2:0];
 reg [31:0] local_size_NO_SHIFT_REG[2:0];
 reg [31:0] work_dim_NO_SHIFT_REG;
 reg [31:0] global_offset_NO_SHIFT_REG[2:0];
 reg [63:0] profile_data_NO_SHIFT_REG;
 reg [31:0] profile_ctrl_NO_SHIFT_REG;
 reg [63:0] profile_start_cycle_NO_SHIFT_REG;
 reg [63:0] profile_stop_cycle_NO_SHIFT_REG;
wire dispatched_all_groups;
wire [31:0] group_id_tmp[2:0];
wire [31:0] global_id_base_out[2:0];
wire start_out;
wire [31:0] local_id[0:0][2:0];
wire [31:0] global_id[0:0][2:0];
wire [31:0] group_id[0:0][2:0];
wire iter_valid_in;
wire iter_stall_out;
wire stall_in;
wire stall_out;
wire valid_in;
wire valid_out;

always @(posedge clock2x or negedge resetn)
begin
	if (~(resetn))
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b0;
	end
	else
	begin
		twoXclock_consumer_NO_SHIFT_REG <= 1'b1;
	end
end



// Work group dispatcher is responsible for issuing work-groups to id iterator(s)
acl_work_group_dispatcher group_dispatcher (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.num_groups(num_groups_NO_SHIFT_REG),
	.local_size(local_size_NO_SHIFT_REG),
	.stall_in(iter_stall_out),
	.valid_out(iter_valid_in),
	.group_id_out(group_id_tmp),
	.global_id_base_out(global_id_base_out),
	.start_out(start_out),
	.dispatched_all_groups(dispatched_all_groups)
);

defparam group_dispatcher.NUM_COPIES = 1;
defparam group_dispatcher.RUN_FOREVER = 0;


// This section of the wrapper implements an Avalon Slave Interface used to configure a kernel invocation.
// The few words words contain the status and the workgroup size registers.
// The remaining addressable space is reserved for kernel arguments.
wire [63:0] bitenable;

assign bitenable[7:0] = (avs_cra_byteenable[0] ? 8'hFF : 8'h0);
assign bitenable[15:8] = (avs_cra_byteenable[1] ? 8'hFF : 8'h0);
assign bitenable[23:16] = (avs_cra_byteenable[2] ? 8'hFF : 8'h0);
assign bitenable[31:24] = (avs_cra_byteenable[3] ? 8'hFF : 8'h0);
assign bitenable[39:32] = (avs_cra_byteenable[4] ? 8'hFF : 8'h0);
assign bitenable[47:40] = (avs_cra_byteenable[5] ? 8'hFF : 8'h0);
assign bitenable[55:48] = (avs_cra_byteenable[6] ? 8'hFF : 8'h0);
assign bitenable[63:56] = (avs_cra_byteenable[7] ? 8'hFF : 8'h0);
assign avs_cra_waitrequest = 1'b0;
assign cra_irq = (status_NO_SHIFT_REG[1] | status_NO_SHIFT_REG[3]);

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		start_NO_SHIFT_REG <= 1'b0;
		started_NO_SHIFT_REG <= 1'b0;
		kernel_arguments_NO_SHIFT_REG <= 448'h0;
		status_NO_SHIFT_REG <= 32'h30000;
		profile_ctrl_NO_SHIFT_REG <= 32'h4;
		profile_start_cycle_NO_SHIFT_REG <= 64'h0;
		profile_stop_cycle_NO_SHIFT_REG <= 64'hFFFFFFFFFFFFFFFF;
		work_dim_NO_SHIFT_REG <= 32'h0;
		workgroup_size_NO_SHIFT_REG <= 32'h0;
		global_size_NO_SHIFT_REG[0] <= 32'h0;
		global_size_NO_SHIFT_REG[1] <= 32'h0;
		global_size_NO_SHIFT_REG[2] <= 32'h0;
		num_groups_NO_SHIFT_REG[0] <= 32'h0;
		num_groups_NO_SHIFT_REG[1] <= 32'h0;
		num_groups_NO_SHIFT_REG[2] <= 32'h0;
		local_size_NO_SHIFT_REG[0] <= 32'h0;
		local_size_NO_SHIFT_REG[1] <= 32'h0;
		local_size_NO_SHIFT_REG[2] <= 32'h0;
		global_offset_NO_SHIFT_REG[0] <= 32'h0;
		global_offset_NO_SHIFT_REG[1] <= 32'h0;
		global_offset_NO_SHIFT_REG[2] <= 32'h0;
	end
	else
	begin
		if (avs_cra_write)
		begin
			case (avs_cra_address)
				5'h0:
				begin
					status_NO_SHIFT_REG[31:16] <= 16'h3;
					status_NO_SHIFT_REG[15:0] <= ((status_NO_SHIFT_REG[15:0] & ~(bitenable[15:0])) | (avs_cra_writedata[15:0] & bitenable[15:0]));
				end

				5'h1:
				begin
					profile_ctrl_NO_SHIFT_REG <= ((profile_ctrl_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h3:
				begin
					profile_start_cycle_NO_SHIFT_REG[31:0] <= ((profile_start_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_start_cycle_NO_SHIFT_REG[63:32] <= ((profile_start_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h4:
				begin
					profile_stop_cycle_NO_SHIFT_REG[31:0] <= ((profile_stop_cycle_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					profile_stop_cycle_NO_SHIFT_REG[63:32] <= ((profile_stop_cycle_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h5:
				begin
					work_dim_NO_SHIFT_REG <= ((work_dim_NO_SHIFT_REG & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					workgroup_size_NO_SHIFT_REG <= ((workgroup_size_NO_SHIFT_REG & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h6:
				begin
					global_size_NO_SHIFT_REG[0] <= ((global_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_size_NO_SHIFT_REG[1] <= ((global_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h7:
				begin
					global_size_NO_SHIFT_REG[2] <= ((global_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[0] <= ((num_groups_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h8:
				begin
					num_groups_NO_SHIFT_REG[1] <= ((num_groups_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					num_groups_NO_SHIFT_REG[2] <= ((num_groups_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h9:
				begin
					local_size_NO_SHIFT_REG[0] <= ((local_size_NO_SHIFT_REG[0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					local_size_NO_SHIFT_REG[1] <= ((local_size_NO_SHIFT_REG[1] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hA:
				begin
					local_size_NO_SHIFT_REG[2] <= ((local_size_NO_SHIFT_REG[2] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[0] <= ((global_offset_NO_SHIFT_REG[0] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hB:
				begin
					global_offset_NO_SHIFT_REG[1] <= ((global_offset_NO_SHIFT_REG[1] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					global_offset_NO_SHIFT_REG[2] <= ((global_offset_NO_SHIFT_REG[2] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hC:
				begin
					kernel_arguments_NO_SHIFT_REG[31:0] <= ((kernel_arguments_NO_SHIFT_REG[31:0] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[63:32] <= ((kernel_arguments_NO_SHIFT_REG[63:32] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hD:
				begin
					kernel_arguments_NO_SHIFT_REG[95:64] <= ((kernel_arguments_NO_SHIFT_REG[95:64] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[127:96] <= ((kernel_arguments_NO_SHIFT_REG[127:96] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hE:
				begin
					kernel_arguments_NO_SHIFT_REG[159:128] <= ((kernel_arguments_NO_SHIFT_REG[159:128] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[191:160] <= ((kernel_arguments_NO_SHIFT_REG[191:160] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'hF:
				begin
					kernel_arguments_NO_SHIFT_REG[223:192] <= ((kernel_arguments_NO_SHIFT_REG[223:192] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[255:224] <= ((kernel_arguments_NO_SHIFT_REG[255:224] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h10:
				begin
					kernel_arguments_NO_SHIFT_REG[287:256] <= ((kernel_arguments_NO_SHIFT_REG[287:256] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[319:288] <= ((kernel_arguments_NO_SHIFT_REG[319:288] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h11:
				begin
					kernel_arguments_NO_SHIFT_REG[351:320] <= ((kernel_arguments_NO_SHIFT_REG[351:320] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[383:352] <= ((kernel_arguments_NO_SHIFT_REG[383:352] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				5'h12:
				begin
					kernel_arguments_NO_SHIFT_REG[415:384] <= ((kernel_arguments_NO_SHIFT_REG[415:384] & ~(bitenable[31:0])) | (avs_cra_writedata[31:0] & bitenable[31:0]));
					kernel_arguments_NO_SHIFT_REG[447:416] <= ((kernel_arguments_NO_SHIFT_REG[447:416] & ~(bitenable[63:32])) | (avs_cra_writedata[63:32] & bitenable[63:32]));
				end

				default:
				begin
				end

			endcase
		end
		else
		begin
			if (status_NO_SHIFT_REG[0])
			begin
				start_NO_SHIFT_REG <= 1'b1;
			end
			if (start_NO_SHIFT_REG)
			begin
				status_NO_SHIFT_REG[0] <= 1'b0;
				started_NO_SHIFT_REG <= 1'b1;
			end
			if (started_NO_SHIFT_REG)
			begin
				start_NO_SHIFT_REG <= 1'b0;
			end
			if (finish)
			begin
				status_NO_SHIFT_REG[1] <= 1'b1;
				started_NO_SHIFT_REG <= 1'b0;
			end
		end
		status_NO_SHIFT_REG[11] <= local_router_hang;
		status_NO_SHIFT_REG[12] <= (|has_a_lsu_active);
		status_NO_SHIFT_REG[13] <= (|has_a_write_pending);
		status_NO_SHIFT_REG[14] <= (|valid_in);
		status_NO_SHIFT_REG[15] <= started_NO_SHIFT_REG;
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		avs_cra_readdata <= 64'h0;
	end
	else
	begin
		case (avs_cra_address)
			5'h0:
			begin
				avs_cra_readdata[31:0] <= status_NO_SHIFT_REG;
				avs_cra_readdata[63:32] <= 32'h0;
			end

			5'h1:
			begin
				avs_cra_readdata[31:0] <= 'x;
				avs_cra_readdata[63:32] <= 32'h0;
			end

			5'h2:
			begin
				avs_cra_readdata[63:0] <= 64'h0;
			end

			5'h3:
			begin
				avs_cra_readdata[63:0] <= 64'h0;
			end

			5'h4:
			begin
				avs_cra_readdata[63:0] <= 64'h0;
			end

			5'h5:
			begin
				avs_cra_readdata[31:0] <= work_dim_NO_SHIFT_REG;
				avs_cra_readdata[63:32] <= workgroup_size_NO_SHIFT_REG;
			end

			5'h6:
			begin
				avs_cra_readdata[31:0] <= global_size_NO_SHIFT_REG[0];
				avs_cra_readdata[63:32] <= global_size_NO_SHIFT_REG[1];
			end

			5'h7:
			begin
				avs_cra_readdata[31:0] <= global_size_NO_SHIFT_REG[2];
				avs_cra_readdata[63:32] <= num_groups_NO_SHIFT_REG[0];
			end

			5'h8:
			begin
				avs_cra_readdata[31:0] <= num_groups_NO_SHIFT_REG[1];
				avs_cra_readdata[63:32] <= num_groups_NO_SHIFT_REG[2];
			end

			5'h9:
			begin
				avs_cra_readdata[31:0] <= local_size_NO_SHIFT_REG[0];
				avs_cra_readdata[63:32] <= local_size_NO_SHIFT_REG[1];
			end

			5'hA:
			begin
				avs_cra_readdata[31:0] <= local_size_NO_SHIFT_REG[2];
				avs_cra_readdata[63:32] <= global_offset_NO_SHIFT_REG[0];
			end

			5'hB:
			begin
				avs_cra_readdata[31:0] <= global_offset_NO_SHIFT_REG[1];
				avs_cra_readdata[63:32] <= global_offset_NO_SHIFT_REG[2];
			end

			5'hC:
			begin
				avs_cra_readdata[31:0] <= kernel_arguments_NO_SHIFT_REG[31:0];
				avs_cra_readdata[63:32] <= kernel_arguments_NO_SHIFT_REG[63:32];
			end

			5'hD:
			begin
				avs_cra_readdata[31:0] <= kernel_arguments_NO_SHIFT_REG[95:64];
				avs_cra_readdata[63:32] <= kernel_arguments_NO_SHIFT_REG[127:96];
			end

			5'hE:
			begin
				avs_cra_readdata[31:0] <= kernel_arguments_NO_SHIFT_REG[159:128];
				avs_cra_readdata[63:32] <= kernel_arguments_NO_SHIFT_REG[191:160];
			end

			5'hF:
			begin
				avs_cra_readdata[31:0] <= kernel_arguments_NO_SHIFT_REG[223:192];
				avs_cra_readdata[63:32] <= kernel_arguments_NO_SHIFT_REG[255:224];
			end

			5'h10:
			begin
				avs_cra_readdata[31:0] <= kernel_arguments_NO_SHIFT_REG[287:256];
				avs_cra_readdata[63:32] <= kernel_arguments_NO_SHIFT_REG[319:288];
			end

			5'h11:
			begin
				avs_cra_readdata[31:0] <= kernel_arguments_NO_SHIFT_REG[351:320];
				avs_cra_readdata[63:32] <= kernel_arguments_NO_SHIFT_REG[383:352];
			end

			5'h12:
			begin
				avs_cra_readdata[31:0] <= kernel_arguments_NO_SHIFT_REG[415:384];
				avs_cra_readdata[63:32] <= kernel_arguments_NO_SHIFT_REG[447:416];
			end

			default:
			begin
				avs_cra_readdata <= status_NO_SHIFT_REG;
			end

		endcase
	end
end

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		avs_cra_readdatavalid <= 1'b0;
	end
	else
	begin
		avs_cra_readdatavalid <= (avs_cra_read & ~(avs_cra_waitrequest));
	end
end


// Handshaking signals used to control data through the pipeline

// Determine when the kernel is finished.
acl_kernel_finish_detector kernel_finish_detector (
	.clock(clock),
	.resetn(resetn),
	.start(start_NO_SHIFT_REG),
	.wg_size(workgroup_size_NO_SHIFT_REG),
	.wg_dispatch_valid_out(iter_valid_in),
	.wg_dispatch_stall_in(iter_stall_out),
	.dispatched_all_groups(dispatched_all_groups),
	.kernel_copy_valid_out(valid_out),
	.kernel_copy_stall_in(stall_in),
	.pending_writes(has_a_write_pending),
	.finish(finish)
);

defparam kernel_finish_detector.NUM_COPIES = 1;
defparam kernel_finish_detector.WG_SIZE_W = 32;

assign stall_in = 1'b0;

// Creating ID iterator and kernel instance for every requested kernel copy

// ID iterator is responsible for iterating over all local ids for given work-groups
acl_id_iterator id_iter_inst0 (
	.clock(clock),
	.resetn(resetn),
	.start(start_out),
	.valid_in(iter_valid_in),
	.stall_out(iter_stall_out),
	.stall_in(stall_out),
	.valid_out(valid_in),
	.group_id_in(group_id_tmp),
	.global_id_base_in(global_id_base_out),
	.local_size(local_size_NO_SHIFT_REG),
	.global_size(global_size_NO_SHIFT_REG),
	.local_id(local_id[0]),
	.global_id(global_id[0]),
	.group_id(group_id[0])
);



// This section instantiates a kernel function block
Matmul_function Matmul_function_inst0 (
	.clock(clock),
	.resetn(resetn),
	.input_global_id_0(global_id[0][0]),
	.input_global_id_1(global_id[0][1]),
	.stall_out(stall_out),
	.valid_in(valid_in),
	.valid_out(valid_out),
	.stall_in(stall_in),
	.workgroup_size(workgroup_size_NO_SHIFT_REG),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_readdata(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_readdata),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_readdatavalid(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_readdatavalid),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_waitrequest(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_waitrequest),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_address(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_address),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_read(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_read),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_write(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_write),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_writeack(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_writeack),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_writedata(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_writedata),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_byteenable(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_byteenable),
	.avm_local_bb2_ld_memcoalesce_m1r_load_0_burstcount(avm_local_bb2_ld_memcoalesce_m1r_load_0_inst0_burstcount),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_readdata(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_readdata),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_readdatavalid(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_readdatavalid),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_waitrequest(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_waitrequest),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_address(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_address),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_read(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_read),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_write(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_write),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_writeack(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_writeack),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_writedata(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_writedata),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_byteenable(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_byteenable),
	.avm_local_bb2_ld_memcoalesce_m1i_load_0_burstcount(avm_local_bb2_ld_memcoalesce_m1i_load_0_inst0_burstcount),
	.avm_local_bb2_ld__readdata(avm_local_bb2_ld__inst0_readdata),
	.avm_local_bb2_ld__readdatavalid(avm_local_bb2_ld__inst0_readdatavalid),
	.avm_local_bb2_ld__waitrequest(avm_local_bb2_ld__inst0_waitrequest),
	.avm_local_bb2_ld__address(avm_local_bb2_ld__inst0_address),
	.avm_local_bb2_ld__read(avm_local_bb2_ld__inst0_read),
	.avm_local_bb2_ld__write(avm_local_bb2_ld__inst0_write),
	.avm_local_bb2_ld__writeack(avm_local_bb2_ld__inst0_writeack),
	.avm_local_bb2_ld__writedata(avm_local_bb2_ld__inst0_writedata),
	.avm_local_bb2_ld__byteenable(avm_local_bb2_ld__inst0_byteenable),
	.avm_local_bb2_ld__burstcount(avm_local_bb2_ld__inst0_burstcount),
	.avm_local_bb2_ld__u1_readdata(avm_local_bb2_ld__u1_inst0_readdata),
	.avm_local_bb2_ld__u1_readdatavalid(avm_local_bb2_ld__u1_inst0_readdatavalid),
	.avm_local_bb2_ld__u1_waitrequest(avm_local_bb2_ld__u1_inst0_waitrequest),
	.avm_local_bb2_ld__u1_address(avm_local_bb2_ld__u1_inst0_address),
	.avm_local_bb2_ld__u1_read(avm_local_bb2_ld__u1_inst0_read),
	.avm_local_bb2_ld__u1_write(avm_local_bb2_ld__u1_inst0_write),
	.avm_local_bb2_ld__u1_writeack(avm_local_bb2_ld__u1_inst0_writeack),
	.avm_local_bb2_ld__u1_writedata(avm_local_bb2_ld__u1_inst0_writedata),
	.avm_local_bb2_ld__u1_byteenable(avm_local_bb2_ld__u1_inst0_byteenable),
	.avm_local_bb2_ld__u1_burstcount(avm_local_bb2_ld__u1_inst0_burstcount),
	.avm_local_bb2_ld__u2_readdata(avm_local_bb2_ld__u2_inst0_readdata),
	.avm_local_bb2_ld__u2_readdatavalid(avm_local_bb2_ld__u2_inst0_readdatavalid),
	.avm_local_bb2_ld__u2_waitrequest(avm_local_bb2_ld__u2_inst0_waitrequest),
	.avm_local_bb2_ld__u2_address(avm_local_bb2_ld__u2_inst0_address),
	.avm_local_bb2_ld__u2_read(avm_local_bb2_ld__u2_inst0_read),
	.avm_local_bb2_ld__u2_write(avm_local_bb2_ld__u2_inst0_write),
	.avm_local_bb2_ld__u2_writeack(avm_local_bb2_ld__u2_inst0_writeack),
	.avm_local_bb2_ld__u2_writedata(avm_local_bb2_ld__u2_inst0_writedata),
	.avm_local_bb2_ld__u2_byteenable(avm_local_bb2_ld__u2_inst0_byteenable),
	.avm_local_bb2_ld__u2_burstcount(avm_local_bb2_ld__u2_inst0_burstcount),
	.avm_local_bb2_ld__u3_readdata(avm_local_bb2_ld__u3_inst0_readdata),
	.avm_local_bb2_ld__u3_readdatavalid(avm_local_bb2_ld__u3_inst0_readdatavalid),
	.avm_local_bb2_ld__u3_waitrequest(avm_local_bb2_ld__u3_inst0_waitrequest),
	.avm_local_bb2_ld__u3_address(avm_local_bb2_ld__u3_inst0_address),
	.avm_local_bb2_ld__u3_read(avm_local_bb2_ld__u3_inst0_read),
	.avm_local_bb2_ld__u3_write(avm_local_bb2_ld__u3_inst0_write),
	.avm_local_bb2_ld__u3_writeack(avm_local_bb2_ld__u3_inst0_writeack),
	.avm_local_bb2_ld__u3_writedata(avm_local_bb2_ld__u3_inst0_writedata),
	.avm_local_bb2_ld__u3_byteenable(avm_local_bb2_ld__u3_inst0_byteenable),
	.avm_local_bb2_ld__u3_burstcount(avm_local_bb2_ld__u3_inst0_burstcount),
	.avm_local_bb3_st_select40_readdata(avm_local_bb3_st_select40_inst0_readdata),
	.avm_local_bb3_st_select40_readdatavalid(avm_local_bb3_st_select40_inst0_readdatavalid),
	.avm_local_bb3_st_select40_waitrequest(avm_local_bb3_st_select40_inst0_waitrequest),
	.avm_local_bb3_st_select40_address(avm_local_bb3_st_select40_inst0_address),
	.avm_local_bb3_st_select40_read(avm_local_bb3_st_select40_inst0_read),
	.avm_local_bb3_st_select40_write(avm_local_bb3_st_select40_inst0_write),
	.avm_local_bb3_st_select40_writeack(avm_local_bb3_st_select40_inst0_writeack),
	.avm_local_bb3_st_select40_writedata(avm_local_bb3_st_select40_inst0_writedata),
	.avm_local_bb3_st_select40_byteenable(avm_local_bb3_st_select40_inst0_byteenable),
	.avm_local_bb3_st_select40_burstcount(avm_local_bb3_st_select40_inst0_burstcount),
	.avm_local_bb3_st_select37_readdata(avm_local_bb3_st_select37_inst0_readdata),
	.avm_local_bb3_st_select37_readdatavalid(avm_local_bb3_st_select37_inst0_readdatavalid),
	.avm_local_bb3_st_select37_waitrequest(avm_local_bb3_st_select37_inst0_waitrequest),
	.avm_local_bb3_st_select37_address(avm_local_bb3_st_select37_inst0_address),
	.avm_local_bb3_st_select37_read(avm_local_bb3_st_select37_inst0_read),
	.avm_local_bb3_st_select37_write(avm_local_bb3_st_select37_inst0_write),
	.avm_local_bb3_st_select37_writeack(avm_local_bb3_st_select37_inst0_writeack),
	.avm_local_bb3_st_select37_writedata(avm_local_bb3_st_select37_inst0_writedata),
	.avm_local_bb3_st_select37_byteenable(avm_local_bb3_st_select37_inst0_byteenable),
	.avm_local_bb3_st_select37_burstcount(avm_local_bb3_st_select37_inst0_burstcount),
	.start(start_out),
	.input_c1f2(kernel_arguments_NO_SHIFT_REG[415:384]),
	.clock2x(clock2x),
	.input_m1r(kernel_arguments_NO_SHIFT_REG[63:0]),
	.input_m1i(kernel_arguments_NO_SHIFT_REG[127:64]),
	.input_col_m2(kernel_arguments_NO_SHIFT_REG[447:416]),
	.input_m2r(kernel_arguments_NO_SHIFT_REG[191:128]),
	.input_m2i(kernel_arguments_NO_SHIFT_REG[255:192]),
	.input_rer(kernel_arguments_NO_SHIFT_REG[319:256]),
	.input_rei(kernel_arguments_NO_SHIFT_REG[383:320]),
	.has_a_write_pending(has_a_write_pending),
	.has_a_lsu_active(has_a_lsu_active)
);



endmodule

//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

module Matmul_sys_cycle_time
	(
		input 		clock,
		input 		resetn,
		output [31:0] 		cur_cycle
	);


 reg [31:0] cur_count_NO_SHIFT_REG;

assign cur_cycle = cur_count_NO_SHIFT_REG;

always @(posedge clock or negedge resetn)
begin
	if (~(resetn))
	begin
		cur_count_NO_SHIFT_REG <= 32'h0;
	end
	else
	begin
		cur_count_NO_SHIFT_REG <= (cur_count_NO_SHIFT_REG + 32'h1);
	end
end

endmodule

